`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 24.01.2020 18:13:04
// Design Name:
// Module Name: test
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////


module simulation();
reg clk,reset;
//reg [5:0]in;
reg [31:0]gamma,row;
wire [63:0]op1,op2;
wire op1_enable;
//wire vaouten;
//integer handle1;
topmod m1 (clk,reset,gamma,row,op1,op2,op1_enable);
/*topmod(clk,reset,gamma,row,op1,op2,op1_enable);*/
initial begin
reset=1;
gamma=0;
row=0;
clk=0;
end

initial
begin
#70 clk=0;
forever #200 clk=~clk;
end

initial begin
#800 reset=0;
end


initial begin
#10000000 $finish;
end

initial
begin 
#450 gamma=32'd1;row=32'd196;
#400 gamma=32'd2;row=32'd157;
#400 gamma=32'd3;row=32'd306;
#400 gamma=32'd3;row=32'd403;
#400 gamma=32'd5;row=32'd174;
#400 gamma=32'd3;row=32'd41;
#400 gamma=32'd4;row=32'd392;
#400 gamma=32'd1;row=32'd292;
#400 gamma=32'd4;row=32'd478;
#400 gamma=32'd2;row=32'd540;
#400 gamma=32'd5;row=32'd416;
#400 gamma=32'd2;row=32'd58;
#400 gamma=32'd4;row=32'd333;
#400 gamma=32'd2;row=32'd241;
#400 gamma=32'd3;row=32'd99;
#400 gamma=32'd1;row=32'd461;
#400 gamma=32'd1;row=32'd196; //jai25
#400 gamma=32'd2;row=32'd157;
#400 gamma=32'd3;row=32'd306;
#400 gamma=32'd3;row=32'd403;
#400 gamma=32'd5;row=32'd174;
#400 gamma=32'd3;row=32'd41;
#400 gamma=32'd4;row=32'd392;
#400 gamma=32'd1;row=32'd292;
#400 gamma=32'd4;row=32'd478;
#400 gamma=32'd2;row=32'd540;
#400 gamma=32'd5;row=32'd416;
#400 gamma=32'd2;row=32'd58;
#400 gamma=32'd4;row=32'd333;
#400 gamma=32'd2;row=32'd241;
#400 gamma=32'd3;row=32'd99;
#400 gamma=32'd1;row=32'd461;
#400 gamma=32'd4;row=32'd297;
#400 gamma=32'd1;row=32'd342;
#400 gamma=32'd5;row=32'd462;
#400 gamma=32'd1;row=32'd194;
#400 gamma=32'd5;row=32'd261;
#400 gamma=32'd5;row=32'd511;
#400 gamma=32'd5;row=32'd233;
#400 gamma=32'd5;row=32'd275;
#400 gamma=32'd2;row=32'd35;
#400 gamma=32'd4;row=32'd381;
#400 gamma=32'd5;row=32'd131;
#400 gamma=32'd2;row=32'd105;
#400 gamma=32'd2;row=32'd193;
#400 gamma=32'd1;row=32'd356;
#400 gamma=32'd5;row=32'd59;
#400 gamma=32'd5;row=32'd307;
#400 gamma=32'd4;row=32'd13;
#400 gamma=32'd2;row=32'd421;
#400 gamma=32'd2;row=32'd331;
#400 gamma=32'd5;row=32'd83;
#400 gamma=32'd2;row=32'd342;
#400 gamma=32'd2;row=32'd243;
#400 gamma=32'd1;row=32'd176;
#400 gamma=32'd5;row=32'd321;
#400 gamma=32'd2;row=32'd493;
#400 gamma=32'd2;row=32'd413;
#400 gamma=32'd1;row=32'd247;
#400 gamma=32'd1;row=32'd326;
#400 gamma=32'd3;row=32'd176;
#400 gamma=32'd3;row=32'd412;
#400 gamma=32'd1;row=32'd337;
#400 gamma=32'd3;row=32'd396;
#400 gamma=32'd5;row=32'd357;
#400 gamma=32'd2;row=32'd375;
#400 gamma=32'd3;row=32'd158;
#400 gamma=32'd5;row=32'd494;
#400 gamma=32'd2;row=32'd438;
#400 gamma=32'd4;row=32'd208;
#400 gamma=32'd1;row=32'd117;
#400 gamma=32'd4;row=32'd505;
#400 gamma=32'd1;row=32'd266;
#400 gamma=32'd1;row=32'd214;
#400 gamma=32'd5;row=32'd347;
#400 gamma=32'd3;row=32'd70;
#400 gamma=32'd5;row=32'd349;
#400 gamma=32'd4;row=32'd170;
#400 gamma=32'd4;row=32'd163;
#400 gamma=32'd5;row=32'd162;
#400 gamma=32'd3;row=32'd460;
#400 gamma=32'd4;row=32'd161;
#400 gamma=32'd1;row=32'd265;
#400 gamma=32'd2;row=32'd499;
#400 gamma=32'd4;row=32'd515;
#400 gamma=32'd2;row=32'd88;
#400 gamma=32'd4;row=32'd150;
#400 gamma=32'd5;row=32'd473;
#400 gamma=32'd4;row=32'd185;
#400 gamma=32'd2;row=32'd30;
#400 gamma=32'd5;row=32'd60;
#400 gamma=32'd1;row=32'd17;
#400 gamma=32'd4;row=32'd475;
#400 gamma=32'd3;row=32'd177;
#400 gamma=32'd1;row=32'd318;
#400 gamma=32'd2;row=32'd450;
#400 gamma=32'd2;row=32'd49;
#400 gamma=32'd2;row=32'd494;
#400 gamma=32'd4;row=32'd215;
#400 gamma=32'd4;row=32'd60;
#400 gamma=32'd2;row=32'd511;
#400 gamma=32'd1;row=32'd318;
#400 gamma=32'd1;row=32'd431;
#400 gamma=32'd2;row=32'd79;
#400 gamma=32'd2;row=32'd137;
#400 gamma=32'd3;row=32'd31;
#400 gamma=32'd2;row=32'd283;
#400 gamma=32'd4;row=32'd451;
#400 gamma=32'd1;row=32'd73;
#400 gamma=32'd2;row=32'd323;
#400 gamma=32'd5;row=32'd259;
#400 gamma=32'd5;row=32'd124;
#400 gamma=32'd4;row=32'd240;
#400 gamma=32'd5;row=32'd409;
#400 gamma=32'd5;row=32'd27;
#400 gamma=32'd5;row=32'd352;
#400 gamma=32'd4;row=32'd526;
#400 gamma=32'd2;row=32'd556;
#400 gamma=32'd1;row=32'd149;
#400 gamma=32'd4;row=32'd446;
#400 gamma=32'd2;row=32'd188;
#400 gamma=32'd4;row=32'd236;
#400 gamma=32'd5;row=32'd104;
#400 gamma=32'd1;row=32'd495;
#400 gamma=32'd3;row=32'd379;
#400 gamma=32'd1;row=32'd272;
#400 gamma=32'd2;row=32'd21;
#400 gamma=32'd1;row=32'd9;
#400 gamma=32'd1;row=32'd397;
#400 gamma=32'd2;row=32'd299;
#400 gamma=32'd3;row=32'd518;
#400 gamma=32'd5;row=32'd266;
#400 gamma=32'd4;row=32'd313;
#400 gamma=32'd2;row=32'd378;
#400 gamma=32'd1;row=32'd173;
#400 gamma=32'd5;row=32'd238;
#400 gamma=32'd2;row=32'd455;
#400 gamma=32'd1;row=32'd70;
#400 gamma=32'd5;row=32'd540;
#400 gamma=32'd2;row=32'd490;
#400 gamma=32'd2;row=32'd31;
#400 gamma=32'd3;row=32'd201;
#400 gamma=32'd5;row=32'd527;
#400 gamma=32'd3;row=32'd425;
#400 gamma=32'd5;row=32'd395;
#400 gamma=32'd5;row=32'd246;
#400 gamma=32'd3;row=32'd306;
#400 gamma=32'd2;row=32'd111;
#400 gamma=32'd3;row=32'd160;
#400 gamma=32'd2;row=32'd146;
#400 gamma=32'd2;row=32'd0;
#400 gamma=32'd5;row=32'd95;
#400 gamma=32'd2;row=32'd373;
#400 gamma=32'd4;row=32'd519;
#400 gamma=32'd1;row=32'd449;
#400 gamma=32'd3;row=32'd429;
#400 gamma=32'd1;row=32'd81;
#400 gamma=32'd2;row=32'd57;
#400 gamma=32'd4;row=32'd512;
#400 gamma=32'd5;row=32'd277;
#400 gamma=32'd2;row=32'd5;
#400 gamma=32'd1;row=32'd125;
#400 gamma=32'd3;row=32'd217;
#400 gamma=32'd1;row=32'd396;
#400 gamma=32'd4;row=32'd452;
#400 gamma=32'd3;row=32'd467;
#400 gamma=32'd3;row=32'd60;
#400 gamma=32'd5;row=32'd161;
#400 gamma=32'd5;row=32'd494;
#400 gamma=32'd1;row=32'd25;
#400 gamma=32'd3;row=32'd374;
#400 gamma=32'd5;row=32'd41;
#400 gamma=32'd1;row=32'd229;
#400 gamma=32'd5;row=32'd123;
#400 gamma=32'd5;row=32'd134;
#400 gamma=32'd2;row=32'd554;
#400 gamma=32'd3;row=32'd138;
#400 gamma=32'd5;row=32'd511;
#400 gamma=32'd3;row=32'd7;
#400 gamma=32'd3;row=32'd207;
#400 gamma=32'd2;row=32'd427;
#400 gamma=32'd4;row=32'd152;
#400 gamma=32'd5;row=32'd280;
#400 gamma=32'd4;row=32'd493;
#400 gamma=32'd5;row=32'd479;
#400 gamma=32'd4;row=32'd430;
#400 gamma=32'd4;row=32'd11;
#400 gamma=32'd3;row=32'd95;
#400 gamma=32'd1;row=32'd487;
#400 gamma=32'd1;row=32'd329;
#400 gamma=32'd2;row=32'd450;
#400 gamma=32'd5;row=32'd129;
#400 gamma=32'd1;row=32'd63;
#400 gamma=32'd2;row=32'd193;
#400 gamma=32'd3;row=32'd281;
#400 gamma=32'd4;row=32'd88;
#400 gamma=32'd1;row=32'd476;
#400 gamma=32'd1;row=32'd291;
#400 gamma=32'd1;row=32'd480;
#400 gamma=32'd4;row=32'd252;
#400 gamma=32'd5;row=32'd353;
#400 gamma=32'd2;row=32'd230;
#400 gamma=32'd1;row=32'd298;
#400 gamma=32'd3;row=32'd500;
#400 gamma=32'd2;row=32'd247;
#400 gamma=32'd3;row=32'd103;
#400 gamma=32'd3;row=32'd91;
#400 gamma=32'd3;row=32'd171;
#400 gamma=32'd2;row=32'd190;
#400 gamma=32'd5;row=32'd359;
#400 gamma=32'd4;row=32'd146;
#400 gamma=32'd1;row=32'd367;
#400 gamma=32'd5;row=32'd1;
#400 gamma=32'd3;row=32'd359;
#400 gamma=32'd5;row=32'd182;
#400 gamma=32'd4;row=32'd231;
#400 gamma=32'd1;row=32'd314;
#400 gamma=32'd3;row=32'd194;
#400 gamma=32'd3;row=32'd304;
#400 gamma=32'd4;row=32'd17;
#400 gamma=32'd1;row=32'd150;
#400 gamma=32'd2;row=32'd189;
#400 gamma=32'd5;row=32'd68;
#400 gamma=32'd3;row=32'd37;
#400 gamma=32'd3;row=32'd480;
#400 gamma=32'd2;row=32'd468;
#400 gamma=32'd4;row=32'd285;
#400 gamma=32'd1;row=32'd288;
#400 gamma=32'd5;row=32'd186;
#400 gamma=32'd1;row=32'd455;
#400 gamma=32'd4;row=32'd206;
#400 gamma=32'd3;row=32'd480;
#400 gamma=32'd2;row=32'd24;
#400 gamma=32'd2;row=32'd29;
#400 gamma=32'd2;row=32'd453;
#400 gamma=32'd1;row=32'd402;
#400 gamma=32'd4;row=32'd356;
#400 gamma=32'd1;row=32'd504;
#400 gamma=32'd3;row=32'd363;
#400 gamma=32'd1;row=32'd150;
#400 gamma=32'd5;row=32'd5;
#400 gamma=32'd4;row=32'd21;
#400 gamma=32'd3;row=32'd268;
#400 gamma=32'd5;row=32'd290;
#400 gamma=32'd4;row=32'd452;
#400 gamma=32'd5;row=32'd472;
#400 gamma=32'd2;row=32'd184;
#400 gamma=32'd3;row=32'd398;
#400 gamma=32'd4;row=32'd211;
#400 gamma=32'd3;row=32'd370;
#400 gamma=32'd2;row=32'd250;
#400 gamma=32'd4;row=32'd496;
#400 gamma=32'd4;row=32'd533;
#400 gamma=32'd3;row=32'd287;
#400 gamma=32'd3;row=32'd127;
#400 gamma=32'd3;row=32'd111;
#400 gamma=32'd2;row=32'd249;
#400 gamma=32'd3;row=32'd273;
#400 gamma=32'd2;row=32'd423;
#400 gamma=32'd5;row=32'd126;
#400 gamma=32'd1;row=32'd87;
#400 gamma=32'd4;row=32'd38;
#400 gamma=32'd2;row=32'd25;
#400 gamma=32'd1;row=32'd75;
#400 gamma=32'd4;row=32'd202;
#400 gamma=32'd2;row=32'd281;
#400 gamma=32'd5;row=32'd210;
#400 gamma=32'd3;row=32'd123;
#400 gamma=32'd3;row=32'd304;
#400 gamma=32'd1;row=32'd290;
#400 gamma=32'd1;row=32'd242;
#400 gamma=32'd4;row=32'd188;
#400 gamma=32'd1;row=32'd85;
#400 gamma=32'd3;row=32'd206;
#400 gamma=32'd4;row=32'd133;
#400 gamma=32'd2;row=32'd284;
#400 gamma=32'd4;row=32'd534;
#400 gamma=32'd4;row=32'd275;
#400 gamma=32'd5;row=32'd366;
#400 gamma=32'd5;row=32'd250;
#400 gamma=32'd3;row=32'd451;
#400 gamma=32'd4;row=32'd53;
#400 gamma=32'd5;row=32'd478;
#400 gamma=32'd2;row=32'd73;
#400 gamma=32'd4;row=32'd127;
#400 gamma=32'd1;row=32'd164;
#400 gamma=32'd5;row=32'd134;
#400 gamma=32'd2;row=32'd332;
#400 gamma=32'd2;row=32'd339;
#400 gamma=32'd4;row=32'd330;
#400 gamma=32'd5;row=32'd12;
#400 gamma=32'd2;row=32'd401;
#400 gamma=32'd4;row=32'd74;
#400 gamma=32'd3;row=32'd523;
#400 gamma=32'd4;row=32'd208;
#400 gamma=32'd5;row=32'd11;
#400 gamma=32'd4;row=32'd449;
#400 gamma=32'd3;row=32'd182;
#400 gamma=32'd3;row=32'd39;
#400 gamma=32'd5;row=32'd447;
#400 gamma=32'd3;row=32'd547;
#400 gamma=32'd5;row=32'd438;
#400 gamma=32'd2;row=32'd33;
#400 gamma=32'd4;row=32'd279;
#400 gamma=32'd5;row=32'd275;
#400 gamma=32'd4;row=32'd10;
#400 gamma=32'd5;row=32'd320;
#400 gamma=32'd5;row=32'd295;
#400 gamma=32'd4;row=32'd448;
#400 gamma=32'd3;row=32'd377;
#400 gamma=32'd3;row=32'd559;
#400 gamma=32'd3;row=32'd366;
#400 gamma=32'd1;row=32'd270;
#400 gamma=32'd5;row=32'd43;
#400 gamma=32'd1;row=32'd420;
#400 gamma=32'd4;row=32'd148;
#400 gamma=32'd4;row=32'd182;
#400 gamma=32'd2;row=32'd368;
#400 gamma=32'd1;row=32'd92;
#400 gamma=32'd4;row=32'd7;
#400 gamma=32'd2;row=32'd467;
#400 gamma=32'd4;row=32'd140;
#400 gamma=32'd5;row=32'd335;
#400 gamma=32'd1;row=32'd113;
#400 gamma=32'd5;row=32'd258;
#400 gamma=32'd1;row=32'd20;
#400 gamma=32'd5;row=32'd263;
#400 gamma=32'd2;row=32'd266;
#400 gamma=32'd4;row=32'd292;
#400 gamma=32'd5;row=32'd135;
#400 gamma=32'd3;row=32'd349;
#400 gamma=32'd5;row=32'd3;
#400 gamma=32'd4;row=32'd224;
#400 gamma=32'd5;row=32'd100;
#400 gamma=32'd2;row=32'd292;
#400 gamma=32'd4;row=32'd261;
#400 gamma=32'd5;row=32'd233;
#400 gamma=32'd1;row=32'd489;
#400 gamma=32'd4;row=32'd269;
#400 gamma=32'd2;row=32'd334;
#400 gamma=32'd3;row=32'd9;
#400 gamma=32'd3;row=32'd544;
#400 gamma=32'd3;row=32'd265;
#400 gamma=32'd2;row=32'd91;
#400 gamma=32'd1;row=32'd368;
#400 gamma=32'd4;row=32'd483;
#400 gamma=32'd4;row=32'd443;
#400 gamma=32'd2;row=32'd11;
#400 gamma=32'd2;row=32'd285;
#400 gamma=32'd1;row=32'd349;
#400 gamma=32'd3;row=32'd336;
#400 gamma=32'd3;row=32'd112;
#400 gamma=32'd5;row=32'd93;
#400 gamma=32'd1;row=32'd134;
#400 gamma=32'd2;row=32'd265;
#400 gamma=32'd2;row=32'd214;
#400 gamma=32'd5;row=32'd275;
#400 gamma=32'd5;row=32'd161;
#400 gamma=32'd4;row=32'd382;
#400 gamma=32'd3;row=32'd389;
#400 gamma=32'd3;row=32'd398;
#400 gamma=32'd5;row=32'd553;
#400 gamma=32'd4;row=32'd471;
#400 gamma=32'd2;row=32'd106;
#400 gamma=32'd2;row=32'd13;
#400 gamma=32'd2;row=32'd55;
#400 gamma=32'd3;row=32'd79;
#400 gamma=32'd3;row=32'd419;
#400 gamma=32'd3;row=32'd530;
#400 gamma=32'd2;row=32'd82;
#400 gamma=32'd1;row=32'd340;
#400 gamma=32'd1;row=32'd224;
#400 gamma=32'd3;row=32'd126;
#400 gamma=32'd1;row=32'd387;
#400 gamma=32'd3;row=32'd423;
#400 gamma=32'd5;row=32'd484;
#400 gamma=32'd2;row=32'd517;
#400 gamma=32'd4;row=32'd212;
#400 gamma=32'd2;row=32'd20;
#400 gamma=32'd5;row=32'd328;
#400 gamma=32'd1;row=32'd18;
#400 gamma=32'd2;row=32'd325;
#400 gamma=32'd3;row=32'd291;
#400 gamma=32'd4;row=32'd290;
#400 gamma=32'd2;row=32'd137;
#400 gamma=32'd1;row=32'd15;
#400 gamma=32'd5;row=32'd374;
#400 gamma=32'd3;row=32'd544;
#400 gamma=32'd5;row=32'd313;
#400 gamma=32'd4;row=32'd370;
#400 gamma=32'd3;row=32'd549;
#400 gamma=32'd2;row=32'd327;
#400 gamma=32'd2;row=32'd193;
#400 gamma=32'd4;row=32'd506;
#400 gamma=32'd1;row=32'd299;
#400 gamma=32'd5;row=32'd73;
#400 gamma=32'd4;row=32'd78;
#400 gamma=32'd3;row=32'd67;
#400 gamma=32'd1;row=32'd366;
#400 gamma=32'd4;row=32'd507;
#400 gamma=32'd4;row=32'd370;
#400 gamma=32'd2;row=32'd27;
#400 gamma=32'd2;row=32'd158;
#400 gamma=32'd1;row=32'd360;
#400 gamma=32'd3;row=32'd58;
#400 gamma=32'd5;row=32'd230;
#400 gamma=32'd2;row=32'd55;
#400 gamma=32'd1;row=32'd221;
#400 gamma=32'd1;row=32'd184;
#400 gamma=32'd4;row=32'd200;
#400 gamma=32'd4;row=32'd339;
#400 gamma=32'd2;row=32'd279;
#400 gamma=32'd3;row=32'd52;
#400 gamma=32'd2;row=32'd89;
#400 gamma=32'd4;row=32'd110;
#400 gamma=32'd2;row=32'd187;
#400 gamma=32'd5;row=32'd102;
#400 gamma=32'd5;row=32'd418;
#400 gamma=32'd1;row=32'd197;
#400 gamma=32'd2;row=32'd336;
#400 gamma=32'd4;row=32'd35;
#400 gamma=32'd2;row=32'd385;
#400 gamma=32'd5;row=32'd508;
#400 gamma=32'd5;row=32'd436;
#400 gamma=32'd1;row=32'd274;
#400 gamma=32'd4;row=32'd209;
#400 gamma=32'd5;row=32'd362;
#400 gamma=32'd3;row=32'd248;
#400 gamma=32'd3;row=32'd357;
#400 gamma=32'd2;row=32'd496;
#400 gamma=32'd4;row=32'd533;
#400 gamma=32'd4;row=32'd221;
#400 gamma=32'd1;row=32'd330;
#400 gamma=32'd4;row=32'd500;
#400 gamma=32'd3;row=32'd497;
#400 gamma=32'd5;row=32'd508;
#400 gamma=32'd2;row=32'd521;
#400 gamma=32'd3;row=32'd196;
#400 gamma=32'd2;row=32'd124;
#400 gamma=32'd3;row=32'd362;
#400 gamma=32'd3;row=32'd350;
#400 gamma=32'd3;row=32'd437;
#400 gamma=32'd3;row=32'd548;
#400 gamma=32'd5;row=32'd456;
#400 gamma=32'd5;row=32'd270;
#400 gamma=32'd2;row=32'd557;
#400 gamma=32'd3;row=32'd45;
#400 gamma=32'd3;row=32'd259;
#400 gamma=32'd3;row=32'd447;
#400 gamma=32'd4;row=32'd83;
#400 gamma=32'd4;row=32'd404;
#400 gamma=32'd2;row=32'd159;
#400 gamma=32'd4;row=32'd434;
#400 gamma=32'd3;row=32'd244;
#400 gamma=32'd2;row=32'd210;
#400 gamma=32'd4;row=32'd18;
#400 gamma=32'd3;row=32'd460;
#400 gamma=32'd5;row=32'd248;
#400 gamma=32'd3;row=32'd441;
#400 gamma=32'd4;row=32'd258;
#400 gamma=32'd5;row=32'd329;
#400 gamma=32'd1;row=32'd264;
#400 gamma=32'd5;row=32'd208;
#400 gamma=32'd1;row=32'd550;
#400 gamma=32'd5;row=32'd427;
#400 gamma=32'd1;row=32'd502;
#400 gamma=32'd5;row=32'd68;
#400 gamma=32'd4;row=32'd302;
#400 gamma=32'd5;row=32'd504;
#400 gamma=32'd5;row=32'd5;
#400 gamma=32'd2;row=32'd419;
#400 gamma=32'd3;row=32'd78;
#400 gamma=32'd2;row=32'd322;
#400 gamma=32'd2;row=32'd76;
#400 gamma=32'd1;row=32'd193;
#400 gamma=32'd4;row=32'd392;
#400 gamma=32'd2;row=32'd395;
#400 gamma=32'd2;row=32'd190;
#400 gamma=32'd2;row=32'd361;
#400 gamma=32'd2;row=32'd432;
#400 gamma=32'd3;row=32'd388;
#400 gamma=32'd1;row=32'd540;
#400 gamma=32'd3;row=32'd112;
#400 gamma=32'd1;row=32'd185;
#400 gamma=32'd3;row=32'd188;
#400 gamma=32'd3;row=32'd454;
#400 gamma=32'd5;row=32'd348;
#400 gamma=32'd2;row=32'd218;
#400 gamma=32'd4;row=32'd195;
#400 gamma=32'd2;row=32'd169;
#400 gamma=32'd1;row=32'd397;
#400 gamma=32'd4;row=32'd300;
#400 gamma=32'd3;row=32'd7;
#400 gamma=32'd3;row=32'd98;
#400 gamma=32'd1;row=32'd274;
#400 gamma=32'd5;row=32'd374;
#400 gamma=32'd5;row=32'd467;
#400 gamma=32'd5;row=32'd304;
#400 gamma=32'd1;row=32'd344;
#400 gamma=32'd3;row=32'd288;
#400 gamma=32'd2;row=32'd537;
#400 gamma=32'd5;row=32'd254;
#400 gamma=32'd4;row=32'd273;
#400 gamma=32'd2;row=32'd145;
#400 gamma=32'd5;row=32'd58;
#400 gamma=32'd1;row=32'd161;
#400 gamma=32'd1;row=32'd70;
#400 gamma=32'd4;row=32'd393;
#400 gamma=32'd3;row=32'd327;
#400 gamma=32'd1;row=32'd239;
#400 gamma=32'd3;row=32'd202;
#400 gamma=32'd5;row=32'd226;
#400 gamma=32'd3;row=32'd487;
#400 gamma=32'd1;row=32'd359;
#400 gamma=32'd3;row=32'd517;
#400 gamma=32'd5;row=32'd459;
#400 gamma=32'd4;row=32'd506;
#400 gamma=32'd4;row=32'd351;
#400 gamma=32'd4;row=32'd465;
#400 gamma=32'd2;row=32'd482;
#400 gamma=32'd4;row=32'd401;
#400 gamma=32'd3;row=32'd293;
#400 gamma=32'd1;row=32'd142;
#400 gamma=32'd5;row=32'd214;
#400 gamma=32'd1;row=32'd406;
#400 gamma=32'd5;row=32'd558;
#400 gamma=32'd4;row=32'd428;
#400 gamma=32'd3;row=32'd508;
#400 gamma=32'd3;row=32'd359;
#400 gamma=32'd3;row=32'd10;
#400 gamma=32'd1;row=32'd455;
#400 gamma=32'd4;row=32'd231;
#400 gamma=32'd2;row=32'd128;
#400 gamma=32'd5;row=32'd510;
#400 gamma=32'd5;row=32'd120;
#400 gamma=32'd1;row=32'd46;
#400 gamma=32'd1;row=32'd541;
#400 gamma=32'd2;row=32'd524;
#400 gamma=32'd2;row=32'd175;
#400 gamma=32'd3;row=32'd128;
#400 gamma=32'd4;row=32'd405;
#400 gamma=32'd3;row=32'd0;
#400 gamma=32'd4;row=32'd313;
#400 gamma=32'd4;row=32'd149;
#400 gamma=32'd2;row=32'd135;
#400 gamma=32'd2;row=32'd324;
#400 gamma=32'd1;row=32'd448;
#400 gamma=32'd1;row=32'd94;
#400 gamma=32'd4;row=32'd5;
#400 gamma=32'd2;row=32'd476;
#400 gamma=32'd3;row=32'd493;
#400 gamma=32'd2;row=32'd130;
#400 gamma=32'd5;row=32'd18;
#400 gamma=32'd1;row=32'd119;
#400 gamma=32'd1;row=32'd115;
#400 gamma=32'd4;row=32'd474;
#400 gamma=32'd3;row=32'd241;
#400 gamma=32'd4;row=32'd288;
#400 gamma=32'd1;row=32'd197;
#400 gamma=32'd5;row=32'd401;
#400 gamma=32'd1;row=32'd140;
#400 gamma=32'd2;row=32'd250;
#400 gamma=32'd3;row=32'd514;
#400 gamma=32'd1;row=32'd457;
#400 gamma=32'd2;row=32'd370;
#400 gamma=32'd3;row=32'd35;
#400 gamma=32'd1;row=32'd84;
#400 gamma=32'd2;row=32'd172;
#400 gamma=32'd4;row=32'd548;
#400 gamma=32'd4;row=32'd544;
#400 gamma=32'd5;row=32'd377;
#400 gamma=32'd2;row=32'd43;
#400 gamma=32'd3;row=32'd92;
#400 gamma=32'd1;row=32'd201;
#400 gamma=32'd2;row=32'd19;
#400 gamma=32'd5;row=32'd237;
#400 gamma=32'd5;row=32'd118;
#400 gamma=32'd1;row=32'd374;
#400 gamma=32'd3;row=32'd82;
#400 gamma=32'd5;row=32'd85;
#400 gamma=32'd1;row=32'd170;
#400 gamma=32'd5;row=32'd183;
#400 gamma=32'd2;row=32'd299;
#400 gamma=32'd3;row=32'd509;
#400 gamma=32'd2;row=32'd79;
#400 gamma=32'd3;row=32'd252;
#400 gamma=32'd3;row=32'd149;
#400 gamma=32'd3;row=32'd408;
#400 gamma=32'd1;row=32'd169;
#400 gamma=32'd3;row=32'd141;
#400 gamma=32'd4;row=32'd190;
#400 gamma=32'd5;row=32'd151;
#400 gamma=32'd5;row=32'd326;
#400 gamma=32'd2;row=32'd361;
#400 gamma=32'd2;row=32'd456;
#400 gamma=32'd4;row=32'd392;
#400 gamma=32'd1;row=32'd328;
#400 gamma=32'd1;row=32'd44;
#400 gamma=32'd3;row=32'd233;
#400 gamma=32'd5;row=32'd189;
#400 gamma=32'd1;row=32'd9;
#400 gamma=32'd5;row=32'd241;
#400 gamma=32'd2;row=32'd473;
#400 gamma=32'd1;row=32'd127;
#400 gamma=32'd4;row=32'd283;
#400 gamma=32'd5;row=32'd131;
#400 gamma=32'd5;row=32'd544;
#400 gamma=32'd1;row=32'd240;
#400 gamma=32'd2;row=32'd12;
#400 gamma=32'd5;row=32'd7;
#400 gamma=32'd1;row=32'd193;
#400 gamma=32'd2;row=32'd439;
#400 gamma=32'd2;row=32'd3;
#400 gamma=32'd4;row=32'd228;
#400 gamma=32'd4;row=32'd78;
#400 gamma=32'd3;row=32'd318;
#400 gamma=32'd1;row=32'd481;
#400 gamma=32'd2;row=32'd312;
#400 gamma=32'd4;row=32'd449;
#400 gamma=32'd5;row=32'd547;
#400 gamma=32'd3;row=32'd379;
#400 gamma=32'd2;row=32'd157;
#400 gamma=32'd1;row=32'd315;
#400 gamma=32'd1;row=32'd148;
#400 gamma=32'd5;row=32'd315;
#400 gamma=32'd4;row=32'd6;
#400 gamma=32'd3;row=32'd498;
#400 gamma=32'd1;row=32'd233;
#400 gamma=32'd2;row=32'd3;
#400 gamma=32'd4;row=32'd224;
#400 gamma=32'd3;row=32'd221;
#400 gamma=32'd3;row=32'd48;
#400 gamma=32'd2;row=32'd204;
#400 gamma=32'd5;row=32'd6;
#400 gamma=32'd1;row=32'd110;
#400 gamma=32'd1;row=32'd225;
#400 gamma=32'd4;row=32'd2;
#400 gamma=32'd4;row=32'd316;
#400 gamma=32'd2;row=32'd281;
#400 gamma=32'd2;row=32'd553;
#400 gamma=32'd3;row=32'd304;
#400 gamma=32'd3;row=32'd296;
#400 gamma=32'd2;row=32'd193;
#400 gamma=32'd1;row=32'd491;
#400 gamma=32'd5;row=32'd382;
#400 gamma=32'd5;row=32'd196;
#400 gamma=32'd3;row=32'd361;
#400 gamma=32'd3;row=32'd370;
#400 gamma=32'd5;row=32'd495;
#400 gamma=32'd1;row=32'd493;
#400 gamma=32'd5;row=32'd172;
#400 gamma=32'd1;row=32'd341;
#400 gamma=32'd5;row=32'd212;
#400 gamma=32'd5;row=32'd527;
#400 gamma=32'd5;row=32'd256;
#400 gamma=32'd4;row=32'd342;
#400 gamma=32'd4;row=32'd86;
#400 gamma=32'd3;row=32'd107;
#400 gamma=32'd1;row=32'd500;
#400 gamma=32'd2;row=32'd328;
#400 gamma=32'd3;row=32'd78;
#400 gamma=32'd4;row=32'd75;
#400 gamma=32'd5;row=32'd166;
#400 gamma=32'd3;row=32'd61;
#400 gamma=32'd4;row=32'd35;
#400 gamma=32'd2;row=32'd506;
#400 gamma=32'd4;row=32'd476;
#400 gamma=32'd5;row=32'd504;
#400 gamma=32'd2;row=32'd181;
#400 gamma=32'd5;row=32'd421;
#400 gamma=32'd1;row=32'd330;
#400 gamma=32'd2;row=32'd344;
#400 gamma=32'd4;row=32'd142;
#400 gamma=32'd3;row=32'd313;
#400 gamma=32'd1;row=32'd371;
#400 gamma=32'd3;row=32'd325;
#400 gamma=32'd4;row=32'd254;
#400 gamma=32'd1;row=32'd98;
#400 gamma=32'd2;row=32'd421;
#400 gamma=32'd5;row=32'd156;
#400 gamma=32'd2;row=32'd345;
#400 gamma=32'd4;row=32'd24;
#400 gamma=32'd3;row=32'd309;
#400 gamma=32'd3;row=32'd126;
#400 gamma=32'd3;row=32'd35;
#400 gamma=32'd5;row=32'd215;
#400 gamma=32'd1;row=32'd482;
#400 gamma=32'd5;row=32'd176;
#400 gamma=32'd4;row=32'd417;
#400 gamma=32'd4;row=32'd184;
#400 gamma=32'd4;row=32'd77;
#400 gamma=32'd4;row=32'd426;
#400 gamma=32'd1;row=32'd161;
#400 gamma=32'd1;row=32'd320;
#400 gamma=32'd3;row=32'd447;
#400 gamma=32'd5;row=32'd395;
#400 gamma=32'd5;row=32'd59;
#400 gamma=32'd5;row=32'd242;
#400 gamma=32'd5;row=32'd501;
#400 gamma=32'd2;row=32'd511;
#400 gamma=32'd3;row=32'd412;
#400 gamma=32'd4;row=32'd369;
#400 gamma=32'd1;row=32'd533;
#400 gamma=32'd2;row=32'd478;
#400 gamma=32'd2;row=32'd75;
#400 gamma=32'd4;row=32'd359;
#400 gamma=32'd1;row=32'd276;
#400 gamma=32'd4;row=32'd427;
#400 gamma=32'd3;row=32'd308;
#400 gamma=32'd5;row=32'd14;
#400 gamma=32'd4;row=32'd251;
#400 gamma=32'd3;row=32'd54;
#400 gamma=32'd3;row=32'd125;
#400 gamma=32'd2;row=32'd296;
#400 gamma=32'd5;row=32'd123;
#400 gamma=32'd1;row=32'd499;
#400 gamma=32'd3;row=32'd451;
#400 gamma=32'd3;row=32'd527;
#400 gamma=32'd5;row=32'd34;
#400 gamma=32'd5;row=32'd110;
#400 gamma=32'd2;row=32'd103;
#400 gamma=32'd3;row=32'd204;
#400 gamma=32'd5;row=32'd87;
#400 gamma=32'd5;row=32'd19;
#400 gamma=32'd5;row=32'd19;
#400 gamma=32'd3;row=32'd396;
#400 gamma=32'd5;row=32'd333;
#400 gamma=32'd4;row=32'd232;
#400 gamma=32'd2;row=32'd1;
#400 gamma=32'd2;row=32'd107;
#400 gamma=32'd3;row=32'd311;
#400 gamma=32'd3;row=32'd236;
#400 gamma=32'd1;row=32'd489;
#400 gamma=32'd5;row=32'd10;
#400 gamma=32'd1;row=32'd209;
#400 gamma=32'd3;row=32'd471;
#400 gamma=32'd1;row=32'd31;
#400 gamma=32'd4;row=32'd549;
#400 gamma=32'd5;row=32'd199;
#400 gamma=32'd4;row=32'd47;
#400 gamma=32'd5;row=32'd215;
#400 gamma=32'd2;row=32'd171;
#400 gamma=32'd2;row=32'd53;
#400 gamma=32'd4;row=32'd159;
#400 gamma=32'd4;row=32'd102;
#400 gamma=32'd1;row=32'd286;
#400 gamma=32'd3;row=32'd14;
#400 gamma=32'd5;row=32'd80;
#400 gamma=32'd2;row=32'd193;
#400 gamma=32'd5;row=32'd382;
#400 gamma=32'd3;row=32'd364;
#400 gamma=32'd4;row=32'd334;
#400 gamma=32'd5;row=32'd194;
#400 gamma=32'd4;row=32'd181;
#400 gamma=32'd4;row=32'd166;
#400 gamma=32'd3;row=32'd2;
#400 gamma=32'd5;row=32'd277;
#400 gamma=32'd2;row=32'd545;
#400 gamma=32'd3;row=32'd550;
#400 gamma=32'd5;row=32'd460;
#400 gamma=32'd4;row=32'd152;
#400 gamma=32'd4;row=32'd402;
#400 gamma=32'd4;row=32'd466;
#400 gamma=32'd3;row=32'd446;
#400 gamma=32'd4;row=32'd134;
#400 gamma=32'd5;row=32'd290;
#400 gamma=32'd5;row=32'd67;
#400 gamma=32'd2;row=32'd386;
#400 gamma=32'd1;row=32'd132;
#400 gamma=32'd4;row=32'd318;
#400 gamma=32'd5;row=32'd517;
#400 gamma=32'd5;row=32'd421;
#400 gamma=32'd4;row=32'd197;
#400 gamma=32'd1;row=32'd224;
#400 gamma=32'd3;row=32'd280;
#400 gamma=32'd5;row=32'd292;
#400 gamma=32'd4;row=32'd78;
#400 gamma=32'd1;row=32'd549;
#400 gamma=32'd1;row=32'd58;
#400 gamma=32'd4;row=32'd176;
#400 gamma=32'd2;row=32'd388;
#400 gamma=32'd2;row=32'd72;
#400 gamma=32'd1;row=32'd133;
#400 gamma=32'd2;row=32'd262;
#400 gamma=32'd5;row=32'd349;
#400 gamma=32'd1;row=32'd510;
#400 gamma=32'd1;row=32'd259;
#400 gamma=32'd2;row=32'd17;
#400 gamma=32'd1;row=32'd473;
#400 gamma=32'd5;row=32'd386;
#400 gamma=32'd4;row=32'd4;
#400 gamma=32'd3;row=32'd478;
#400 gamma=32'd2;row=32'd456;
#400 gamma=32'd4;row=32'd257;
#400 gamma=32'd3;row=32'd444;
#400 gamma=32'd4;row=32'd489;
#400 gamma=32'd3;row=32'd456;
#400 gamma=32'd5;row=32'd417;
#400 gamma=32'd4;row=32'd277;
#400 gamma=32'd3;row=32'd41;
#400 gamma=32'd5;row=32'd50;
#400 gamma=32'd4;row=32'd220;
#400 gamma=32'd2;row=32'd493;
#400 gamma=32'd2;row=32'd296;
#400 gamma=32'd4;row=32'd357;
#400 gamma=32'd2;row=32'd304;
#400 gamma=32'd1;row=32'd249;
#400 gamma=32'd4;row=32'd329;
#400 gamma=32'd4;row=32'd402;
#400 gamma=32'd4;row=32'd381;
#400 gamma=32'd2;row=32'd298;
#400 gamma=32'd1;row=32'd196;
#400 gamma=32'd1;row=32'd158;
#400 gamma=32'd4;row=32'd529;
#400 gamma=32'd3;row=32'd174;
#400 gamma=32'd2;row=32'd461;
#400 gamma=32'd5;row=32'd198;
#400 gamma=32'd4;row=32'd458;
#400 gamma=32'd4;row=32'd51;
#400 gamma=32'd5;row=32'd295;
#400 gamma=32'd5;row=32'd341;
#400 gamma=32'd2;row=32'd179;
#400 gamma=32'd3;row=32'd127;
#400 gamma=32'd4;row=32'd432;
#400 gamma=32'd4;row=32'd505;
#400 gamma=32'd5;row=32'd317;
#400 gamma=32'd1;row=32'd106;
#400 gamma=32'd5;row=32'd365;
#400 gamma=32'd2;row=32'd215;
#400 gamma=32'd5;row=32'd548;
#400 gamma=32'd4;row=32'd333;
#400 gamma=32'd1;row=32'd7;
#400 gamma=32'd3;row=32'd35;
#400 gamma=32'd1;row=32'd201;
#400 gamma=32'd5;row=32'd99;
#400 gamma=32'd4;row=32'd146;
#400 gamma=32'd5;row=32'd500;
#400 gamma=32'd1;row=32'd47;
#400 gamma=32'd5;row=32'd405;
#400 gamma=32'd4;row=32'd447;
#400 gamma=32'd1;row=32'd347;
#400 gamma=32'd3;row=32'd535;
#400 gamma=32'd4;row=32'd445;
#400 gamma=32'd1;row=32'd169;
#400 gamma=32'd4;row=32'd261;
#400 gamma=32'd1;row=32'd376;
#400 gamma=32'd4;row=32'd346;
#400 gamma=32'd5;row=32'd252;
#400 gamma=32'd2;row=32'd191;
#400 gamma=32'd2;row=32'd506;
#400 gamma=32'd3;row=32'd555;
#400 gamma=32'd2;row=32'd548;
#400 gamma=32'd4;row=32'd389;
#400 gamma=32'd4;row=32'd512;
#400 gamma=32'd1;row=32'd381;
#400 gamma=32'd3;row=32'd170;
#400 gamma=32'd2;row=32'd110;
#400 gamma=32'd4;row=32'd347;
#400 gamma=32'd2;row=32'd284;
#400 gamma=32'd1;row=32'd79;
#400 gamma=32'd2;row=32'd523;
#400 gamma=32'd3;row=32'd243;
#400 gamma=32'd2;row=32'd470;
#400 gamma=32'd3;row=32'd366;
#400 gamma=32'd1;row=32'd438;
#400 gamma=32'd2;row=32'd559;
#400 gamma=32'd4;row=32'd488;
#400 gamma=32'd5;row=32'd264;
#400 gamma=32'd2;row=32'd501;
#400 gamma=32'd1;row=32'd435;
#400 gamma=32'd3;row=32'd58;
#400 gamma=32'd3;row=32'd194;
#400 gamma=32'd5;row=32'd526;
#400 gamma=32'd3;row=32'd42;
#400 gamma=32'd2;row=32'd317;
#400 gamma=32'd4;row=32'd551;
#400 gamma=32'd5;row=32'd54;
#400 gamma=32'd2;row=32'd321;
#400 gamma=32'd5;row=32'd536;
#400 gamma=32'd2;row=32'd262;
#400 gamma=32'd3;row=32'd365;
#400 gamma=32'd2;row=32'd334;
#400 gamma=32'd3;row=32'd541;
#400 gamma=32'd4;row=32'd138;
#400 gamma=32'd2;row=32'd8;
#400 gamma=32'd1;row=32'd120;
#400 gamma=32'd1;row=32'd57;
#400 gamma=32'd5;row=32'd344;
#400 gamma=32'd5;row=32'd253;
#400 gamma=32'd5;row=32'd515;
#400 gamma=32'd4;row=32'd325;
#400 gamma=32'd5;row=32'd240;
#400 gamma=32'd4;row=32'd421;
#400 gamma=32'd4;row=32'd494;
#400 gamma=32'd3;row=32'd411;
#400 gamma=32'd1;row=32'd178;
#400 gamma=32'd4;row=32'd481;
#400 gamma=32'd3;row=32'd90;
#400 gamma=32'd3;row=32'd553;
#400 gamma=32'd4;row=32'd430;
#400 gamma=32'd2;row=32'd259;
#400 gamma=32'd5;row=32'd468;
#400 gamma=32'd5;row=32'd204;
#400 gamma=32'd2;row=32'd485;
#400 gamma=32'd1;row=32'd122;
#400 gamma=32'd2;row=32'd167;
#400 gamma=32'd4;row=32'd389;
#400 gamma=32'd5;row=32'd50;
#400 gamma=32'd1;row=32'd192;
#400 gamma=32'd3;row=32'd169;
#400 gamma=32'd4;row=32'd352;
#400 gamma=32'd1;row=32'd31;
#400 gamma=32'd3;row=32'd156;
#400 gamma=32'd3;row=32'd538;
#400 gamma=32'd5;row=32'd417;
#400 gamma=32'd5;row=32'd425;
#400 gamma=32'd1;row=32'd283;
#400 gamma=32'd5;row=32'd23;
#400 gamma=32'd4;row=32'd19;
#400 gamma=32'd1;row=32'd414;
#400 gamma=32'd4;row=32'd194;
#400 gamma=32'd1;row=32'd282;
#400 gamma=32'd5;row=32'd178;
#400 gamma=32'd5;row=32'd4;
#400 gamma=32'd1;row=32'd44;
#400 gamma=32'd3;row=32'd312;
#400 gamma=32'd4;row=32'd51;
#400 gamma=32'd1;row=32'd481;
#400 gamma=32'd3;row=32'd44;
#400 gamma=32'd1;row=32'd429;
#400 gamma=32'd5;row=32'd58;
#400 gamma=32'd5;row=32'd273;
#400 gamma=32'd2;row=32'd492;
#400 gamma=32'd1;row=32'd163;
#400 gamma=32'd3;row=32'd553;
#400 gamma=32'd5;row=32'd356;
#400 gamma=32'd3;row=32'd233;
#400 gamma=32'd4;row=32'd339;
#400 gamma=32'd3;row=32'd96;
#400 gamma=32'd4;row=32'd118;
#400 gamma=32'd3;row=32'd234;
#400 gamma=32'd1;row=32'd301;
#400 gamma=32'd2;row=32'd215;
#400 gamma=32'd1;row=32'd500;
#400 gamma=32'd3;row=32'd487;
#400 gamma=32'd2;row=32'd461;
#400 gamma=32'd1;row=32'd122;
#400 gamma=32'd5;row=32'd59;
#400 gamma=32'd3;row=32'd111;
#400 gamma=32'd2;row=32'd151;
#400 gamma=32'd1;row=32'd474;
#400 gamma=32'd3;row=32'd18;
#400 gamma=32'd4;row=32'd331;
#400 gamma=32'd3;row=32'd459;
#400 gamma=32'd4;row=32'd441;
#400 gamma=32'd1;row=32'd428;
#400 gamma=32'd5;row=32'd300;
#400 gamma=32'd4;row=32'd282;
#400 gamma=32'd5;row=32'd398;
#400 gamma=32'd5;row=32'd416;
#400 gamma=32'd1;row=32'd218;
#400 gamma=32'd4;row=32'd319;
#400 gamma=32'd2;row=32'd83;
#400 gamma=32'd1;row=32'd451;
#400 gamma=32'd5;row=32'd418;
#400 gamma=32'd2;row=32'd466;
#400 gamma=32'd4;row=32'd11;
#400 gamma=32'd5;row=32'd3;
#400 gamma=32'd4;row=32'd552;
#400 gamma=32'd5;row=32'd534;
#400 gamma=32'd4;row=32'd309;
#400 gamma=32'd1;row=32'd69;
#400 gamma=32'd2;row=32'd466;
#400 gamma=32'd2;row=32'd165;
#400 gamma=32'd4;row=32'd370;
#400 gamma=32'd2;row=32'd467;
#400 gamma=32'd5;row=32'd117;
#400 gamma=32'd1;row=32'd485;
#400 gamma=32'd2;row=32'd34;
#400 gamma=32'd2;row=32'd140;
#400 gamma=32'd4;row=32'd288;
#400 gamma=32'd4;row=32'd456;
#400 gamma=32'd5;row=32'd210;
#400 gamma=32'd5;row=32'd173;
#400 gamma=32'd3;row=32'd389;
#400 gamma=32'd4;row=32'd378;
#400 gamma=32'd1;row=32'd66;
#400 gamma=32'd5;row=32'd219;
#400 gamma=32'd1;row=32'd175;
#400 gamma=32'd5;row=32'd549;
#400 gamma=32'd5;row=32'd107;
#400 gamma=32'd2;row=32'd451;
#400 gamma=32'd3;row=32'd4;
#400 gamma=32'd2;row=32'd535;
#400 gamma=32'd5;row=32'd201;
#400 gamma=32'd3;row=32'd434;
#400 gamma=32'd4;row=32'd278;
#400 gamma=32'd3;row=32'd468;
#400 gamma=32'd3;row=32'd547;
#400 gamma=32'd5;row=32'd24;
#400 gamma=32'd5;row=32'd487;
#400 gamma=32'd2;row=32'd366;
#400 gamma=32'd1;row=32'd251;
#400 gamma=32'd3;row=32'd491;
#400 gamma=32'd2;row=32'd510;
#400 gamma=32'd4;row=32'd526;
#400 gamma=32'd2;row=32'd503;
#400 gamma=32'd1;row=32'd101;
#400 gamma=32'd5;row=32'd16;
#400 gamma=32'd3;row=32'd251;
#400 gamma=32'd1;row=32'd166;
#400 gamma=32'd1;row=32'd423;
#400 gamma=32'd1;row=32'd35;
#400 gamma=32'd3;row=32'd238;
#400 gamma=32'd2;row=32'd211;
#400 gamma=32'd1;row=32'd499;
#400 gamma=32'd3;row=32'd39;
#400 gamma=32'd1;row=32'd276;
#400 gamma=32'd2;row=32'd450;
#400 gamma=32'd1;row=32'd171;
#400 gamma=32'd3;row=32'd20;
#400 gamma=32'd3;row=32'd144;
#400 gamma=32'd4;row=32'd145;
#400 gamma=32'd2;row=32'd150;
#400 gamma=32'd1;row=32'd419;
#400 gamma=32'd4;row=32'd201;
#400 gamma=32'd3;row=32'd107;
#400 gamma=32'd4;row=32'd541;
#400 gamma=32'd3;row=32'd322;
#400 gamma=32'd2;row=32'd307;
#400 gamma=32'd1;row=32'd503;
#400 gamma=32'd2;row=32'd354;
#400 gamma=32'd1;row=32'd390;
#400 gamma=32'd4;row=32'd498;
#400 gamma=32'd1;row=32'd241;
#400 gamma=32'd5;row=32'd509;
#400 gamma=32'd4;row=32'd213;
#400 gamma=32'd5;row=32'd553;
#400 gamma=32'd2;row=32'd291;
#400 gamma=32'd3;row=32'd382;
#400 gamma=32'd2;row=32'd333;
#400 gamma=32'd1;row=32'd187;
#400 gamma=32'd1;row=32'd226;
#400 gamma=32'd5;row=32'd320;
#400 gamma=32'd5;row=32'd92;
#400 gamma=32'd2;row=32'd62;
#400 gamma=32'd2;row=32'd513;
#400 gamma=32'd5;row=32'd48;
#400 gamma=32'd3;row=32'd412;
#400 gamma=32'd5;row=32'd267;
#400 gamma=32'd2;row=32'd279;
#400 gamma=32'd1;row=32'd217;
#400 gamma=32'd5;row=32'd2;
#400 gamma=32'd2;row=32'd155;
#400 gamma=32'd2;row=32'd546;
#400 gamma=32'd3;row=32'd466;
#400 gamma=32'd2;row=32'd363;
#400 gamma=32'd4;row=32'd94;
#400 gamma=32'd4;row=32'd116;
#400 gamma=32'd1;row=32'd210;
#400 gamma=32'd4;row=32'd61;
#400 gamma=32'd3;row=32'd94;
#400 gamma=32'd5;row=32'd87;
#400 gamma=32'd1;row=32'd449;
#400 gamma=32'd1;row=32'd310;
#400 gamma=32'd3;row=32'd319;
#400 gamma=32'd3;row=32'd130;
#400 gamma=32'd4;row=32'd140;
#400 gamma=32'd2;row=32'd200;
#400 gamma=32'd3;row=32'd107;
#400 gamma=32'd2;row=32'd177;
#400 gamma=32'd3;row=32'd456;
#400 gamma=32'd5;row=32'd521;
#400 gamma=32'd5;row=32'd496;
#400 gamma=32'd2;row=32'd159;
#400 gamma=32'd4;row=32'd450;
#400 gamma=32'd3;row=32'd390;
#400 gamma=32'd3;row=32'd381;
#400 gamma=32'd1;row=32'd525;
#400 gamma=32'd5;row=32'd477;
#400 gamma=32'd5;row=32'd215;
#400 gamma=32'd1;row=32'd157;
#400 gamma=32'd3;row=32'd492;
#400 gamma=32'd4;row=32'd328;
#400 gamma=32'd4;row=32'd432;
#400 gamma=32'd2;row=32'd72;
#400 gamma=32'd1;row=32'd104;
#400 gamma=32'd2;row=32'd470;
#400 gamma=32'd3;row=32'd449;
#400 gamma=32'd4;row=32'd489;
#400 gamma=32'd5;row=32'd65;
#400 gamma=32'd5;row=32'd206;
#400 gamma=32'd4;row=32'd376;
#400 gamma=32'd1;row=32'd505;
#400 gamma=32'd1;row=32'd213;
#400 gamma=32'd1;row=32'd8;
#400 gamma=32'd4;row=32'd58;
#400 gamma=32'd3;row=32'd229;
#400 gamma=32'd2;row=32'd525;
#400 gamma=32'd1;row=32'd279;
#400 gamma=32'd2;row=32'd62;
#400 gamma=32'd4;row=32'd147;
#400 gamma=32'd5;row=32'd299;
#400 gamma=32'd5;row=32'd40;
#400 gamma=32'd1;row=32'd513;
#400 gamma=32'd5;row=32'd440;
#400 gamma=32'd5;row=32'd469;
#400 gamma=32'd2;row=32'd398;
#400 gamma=32'd3;row=32'd65;
#400 gamma=32'd2;row=32'd195;
#400 gamma=32'd2;row=32'd38;
#400 gamma=32'd2;row=32'd2;
#400 gamma=32'd4;row=32'd452;
#400 gamma=32'd5;row=32'd84;
#400 gamma=32'd3;row=32'd127;
#400 gamma=32'd4;row=32'd491;
#400 gamma=32'd3;row=32'd321;
#400 gamma=32'd1;row=32'd389;
#400 gamma=32'd4;row=32'd273;
#400 gamma=32'd3;row=32'd196;
#400 gamma=32'd4;row=32'd252;
#400 gamma=32'd4;row=32'd204;
#400 gamma=32'd3;row=32'd42;
#400 gamma=32'd3;row=32'd550;
#400 gamma=32'd5;row=32'd503;
#400 gamma=32'd3;row=32'd65;
#400 gamma=32'd2;row=32'd402;
#400 gamma=32'd3;row=32'd482;
#400 gamma=32'd2;row=32'd11;
#400 gamma=32'd4;row=32'd97;
#400 gamma=32'd1;row=32'd499;
#400 gamma=32'd2;row=32'd26;
#400 gamma=32'd3;row=32'd207;
#400 gamma=32'd2;row=32'd154;
#400 gamma=32'd1;row=32'd536;
#400 gamma=32'd1;row=32'd504;
#400 gamma=32'd1;row=32'd101;
#400 gamma=32'd4;row=32'd71;
#400 gamma=32'd4;row=32'd76;
#400 gamma=32'd4;row=32'd437;
#400 gamma=32'd3;row=32'd166;
#400 gamma=32'd4;row=32'd170;
#400 gamma=32'd1;row=32'd501;
#400 gamma=32'd3;row=32'd546;
#400 gamma=32'd3;row=32'd83;
#400 gamma=32'd1;row=32'd49;
#400 gamma=32'd3;row=32'd251;
#400 gamma=32'd1;row=32'd4;
#400 gamma=32'd4;row=32'd71;
#400 gamma=32'd2;row=32'd525;
#400 gamma=32'd4;row=32'd451;
#400 gamma=32'd4;row=32'd298;
#400 gamma=32'd2;row=32'd210;
#400 gamma=32'd2;row=32'd548;
#400 gamma=32'd3;row=32'd421;
#400 gamma=32'd3;row=32'd220;
#400 gamma=32'd5;row=32'd410;
#400 gamma=32'd1;row=32'd48;
#400 gamma=32'd2;row=32'd443;
#400 gamma=32'd3;row=32'd352;
#400 gamma=32'd2;row=32'd131;
#400 gamma=32'd5;row=32'd430;
#400 gamma=32'd3;row=32'd106;
#400 gamma=32'd5;row=32'd385;
#400 gamma=32'd2;row=32'd357;
#400 gamma=32'd2;row=32'd542;
#400 gamma=32'd1;row=32'd291;
#400 gamma=32'd5;row=32'd490;
#400 gamma=32'd4;row=32'd56;
#400 gamma=32'd1;row=32'd411;
#400 gamma=32'd3;row=32'd74;
#400 gamma=32'd5;row=32'd189;
#400 gamma=32'd3;row=32'd551;
#400 gamma=32'd2;row=32'd205;
#400 gamma=32'd3;row=32'd300;
#400 gamma=32'd3;row=32'd236;
#400 gamma=32'd1;row=32'd254;
#400 gamma=32'd4;row=32'd215;
#400 gamma=32'd4;row=32'd488;
#400 gamma=32'd4;row=32'd38;
#400 gamma=32'd4;row=32'd29;
#400 gamma=32'd4;row=32'd554;
#400 gamma=32'd4;row=32'd119;
#400 gamma=32'd4;row=32'd183;
#400 gamma=32'd5;row=32'd467;
#400 gamma=32'd1;row=32'd172;
#400 gamma=32'd4;row=32'd212;
#400 gamma=32'd2;row=32'd528;
#400 gamma=32'd1;row=32'd73;
#400 gamma=32'd5;row=32'd353;
#400 gamma=32'd1;row=32'd332;
#400 gamma=32'd2;row=32'd401;
#400 gamma=32'd1;row=32'd219;
#400 gamma=32'd4;row=32'd259;
#400 gamma=32'd2;row=32'd479;
#400 gamma=32'd1;row=32'd220;
#400 gamma=32'd3;row=32'd62;
#400 gamma=32'd1;row=32'd339;
#400 gamma=32'd1;row=32'd146;
#400 gamma=32'd1;row=32'd317;
#400 gamma=32'd4;row=32'd66;
#400 gamma=32'd1;row=32'd512;
#400 gamma=32'd4;row=32'd395;
#400 gamma=32'd4;row=32'd244;
#400 gamma=32'd3;row=32'd178;
#400 gamma=32'd5;row=32'd443;
#400 gamma=32'd4;row=32'd279;
#400 gamma=32'd5;row=32'd484;
#400 gamma=32'd3;row=32'd158;
#400 gamma=32'd2;row=32'd542;
#400 gamma=32'd5;row=32'd506;
#400 gamma=32'd4;row=32'd472;
#400 gamma=32'd1;row=32'd365;
#400 gamma=32'd5;row=32'd435;
#400 gamma=32'd1;row=32'd310;
#400 gamma=32'd3;row=32'd399;
#400 gamma=32'd2;row=32'd301;
#400 gamma=32'd5;row=32'd443;
#400 gamma=32'd2;row=32'd418;
#400 gamma=32'd4;row=32'd222;
#400 gamma=32'd3;row=32'd161;
#400 gamma=32'd1;row=32'd259;
#400 gamma=32'd4;row=32'd390;
#400 gamma=32'd1;row=32'd227;
#400 gamma=32'd2;row=32'd128;
#400 gamma=32'd1;row=32'd28;
#400 gamma=32'd5;row=32'd98;
#400 gamma=32'd4;row=32'd219;
#400 gamma=32'd3;row=32'd547;
#400 gamma=32'd5;row=32'd479;
#400 gamma=32'd1;row=32'd492;
#400 gamma=32'd3;row=32'd420;
#400 gamma=32'd4;row=32'd466;
#400 gamma=32'd1;row=32'd20;
#400 gamma=32'd4;row=32'd101;
#400 gamma=32'd5;row=32'd47;
#400 gamma=32'd3;row=32'd145;
#400 gamma=32'd1;row=32'd245;
#400 gamma=32'd3;row=32'd540;
#400 gamma=32'd3;row=32'd102;
#400 gamma=32'd3;row=32'd455;
#400 gamma=32'd4;row=32'd537;
#400 gamma=32'd2;row=32'd357;
#400 gamma=32'd1;row=32'd188;
#400 gamma=32'd5;row=32'd41;
#400 gamma=32'd4;row=32'd20;
#400 gamma=32'd5;row=32'd505;
#400 gamma=32'd1;row=32'd6;
#400 gamma=32'd2;row=32'd317;
#400 gamma=32'd2;row=32'd519;
#400 gamma=32'd2;row=32'd57;
#400 gamma=32'd1;row=32'd536;
#400 gamma=32'd1;row=32'd339;
#400 gamma=32'd1;row=32'd100;
#400 gamma=32'd4;row=32'd83;
#400 gamma=32'd4;row=32'd407;
#400 gamma=32'd2;row=32'd519;
#400 gamma=32'd2;row=32'd23;
#400 gamma=32'd1;row=32'd439;
#400 gamma=32'd3;row=32'd442;
#400 gamma=32'd2;row=32'd179;
#400 gamma=32'd2;row=32'd371;
#400 gamma=32'd4;row=32'd277;
#400 gamma=32'd4;row=32'd334;
#400 gamma=32'd4;row=32'd422;
#400 gamma=32'd5;row=32'd85;
#400 gamma=32'd1;row=32'd510;
#400 gamma=32'd1;row=32'd441;
#400 gamma=32'd1;row=32'd259;
#400 gamma=32'd3;row=32'd5;
#400 gamma=32'd5;row=32'd220;
#400 gamma=32'd2;row=32'd351;
#400 gamma=32'd1;row=32'd172;
#400 gamma=32'd3;row=32'd109;
#400 gamma=32'd2;row=32'd500;
#400 gamma=32'd2;row=32'd0;
#400 gamma=32'd3;row=32'd278;
#400 gamma=32'd3;row=32'd215;
#400 gamma=32'd3;row=32'd69;
#400 gamma=32'd4;row=32'd122;
#400 gamma=32'd3;row=32'd470;
#400 gamma=32'd2;row=32'd481;
#400 gamma=32'd2;row=32'd507;
#400 gamma=32'd1;row=32'd308;
#400 gamma=32'd5;row=32'd299;
#400 gamma=32'd3;row=32'd280;
#400 gamma=32'd1;row=32'd270;
#400 gamma=32'd1;row=32'd337;
#400 gamma=32'd3;row=32'd78;
#400 gamma=32'd5;row=32'd344;
#400 gamma=32'd5;row=32'd40;
#400 gamma=32'd3;row=32'd351;
#400 gamma=32'd2;row=32'd151;
#400 gamma=32'd5;row=32'd422;
#400 gamma=32'd3;row=32'd59;
#400 gamma=32'd3;row=32'd488;
#400 gamma=32'd2;row=32'd450;
#400 gamma=32'd4;row=32'd100;
#400 gamma=32'd2;row=32'd85;
#400 gamma=32'd5;row=32'd100;
#400 gamma=32'd1;row=32'd262;
#400 gamma=32'd2;row=32'd313;
#400 gamma=32'd2;row=32'd450;
#400 gamma=32'd3;row=32'd117;
#400 gamma=32'd3;row=32'd273;
#400 gamma=32'd5;row=32'd537;
#400 gamma=32'd3;row=32'd167;
#400 gamma=32'd5;row=32'd51;
#400 gamma=32'd3;row=32'd539;
#400 gamma=32'd4;row=32'd24;
#400 gamma=32'd4;row=32'd314;
#400 gamma=32'd4;row=32'd22;
#400 gamma=32'd1;row=32'd25;
#400 gamma=32'd1;row=32'd439;
#400 gamma=32'd3;row=32'd257;
#400 gamma=32'd3;row=32'd73;
#400 gamma=32'd3;row=32'd283;
#400 gamma=32'd1;row=32'd357;
#400 gamma=32'd1;row=32'd81;
#400 gamma=32'd3;row=32'd485;
#400 gamma=32'd4;row=32'd117;
#400 gamma=32'd4;row=32'd227;
#400 gamma=32'd5;row=32'd394;
#400 gamma=32'd4;row=32'd263;
#400 gamma=32'd1;row=32'd160;
#400 gamma=32'd2;row=32'd528;
#400 gamma=32'd5;row=32'd39;
#400 gamma=32'd1;row=32'd489;
#400 gamma=32'd5;row=32'd112;
#400 gamma=32'd1;row=32'd284;
#400 gamma=32'd2;row=32'd120;
#400 gamma=32'd2;row=32'd495;
#400 gamma=32'd1;row=32'd67;
#400 gamma=32'd2;row=32'd114;
#400 gamma=32'd1;row=32'd510;
#400 gamma=32'd2;row=32'd98;
#400 gamma=32'd1;row=32'd511;
#400 gamma=32'd3;row=32'd48;
#400 gamma=32'd4;row=32'd165;
#400 gamma=32'd4;row=32'd545;
#400 gamma=32'd3;row=32'd153;
#400 gamma=32'd5;row=32'd211;
#400 gamma=32'd2;row=32'd167;
#400 gamma=32'd5;row=32'd497;
#400 gamma=32'd4;row=32'd91;
#400 gamma=32'd5;row=32'd133;
#400 gamma=32'd3;row=32'd94;
#400 gamma=32'd1;row=32'd160;
#400 gamma=32'd5;row=32'd251;
#400 gamma=32'd3;row=32'd92;
#400 gamma=32'd5;row=32'd554;
#400 gamma=32'd1;row=32'd546;
#400 gamma=32'd4;row=32'd470;
#400 gamma=32'd4;row=32'd487;
#400 gamma=32'd5;row=32'd448;
#400 gamma=32'd3;row=32'd475;
#400 gamma=32'd4;row=32'd134;
#400 gamma=32'd1;row=32'd534;
#400 gamma=32'd3;row=32'd227;
#400 gamma=32'd3;row=32'd84;
#400 gamma=32'd1;row=32'd88;
#400 gamma=32'd2;row=32'd366;
#400 gamma=32'd3;row=32'd368;
#400 gamma=32'd3;row=32'd2;
#400 gamma=32'd1;row=32'd485;
#400 gamma=32'd3;row=32'd231;
#400 gamma=32'd5;row=32'd452;
#400 gamma=32'd3;row=32'd12;
#400 gamma=32'd1;row=32'd8;
#400 gamma=32'd1;row=32'd505;
#400 gamma=32'd1;row=32'd193;
#400 gamma=32'd4;row=32'd107;
#400 gamma=32'd1;row=32'd520;
#400 gamma=32'd1;row=32'd532;
#400 gamma=32'd4;row=32'd49;
#400 gamma=32'd1;row=32'd467;
#400 gamma=32'd1;row=32'd513;
#400 gamma=32'd3;row=32'd233;
#400 gamma=32'd1;row=32'd505;
#400 gamma=32'd3;row=32'd63;
#400 gamma=32'd4;row=32'd235;
#400 gamma=32'd3;row=32'd7;
#400 gamma=32'd3;row=32'd259;
#400 gamma=32'd5;row=32'd273;
#400 gamma=32'd4;row=32'd454;
#400 gamma=32'd3;row=32'd105;
#400 gamma=32'd1;row=32'd353;
#400 gamma=32'd2;row=32'd28;
#400 gamma=32'd1;row=32'd85;
#400 gamma=32'd1;row=32'd191;
#400 gamma=32'd4;row=32'd255;
#400 gamma=32'd2;row=32'd299;
#400 gamma=32'd4;row=32'd540;
#400 gamma=32'd5;row=32'd134;
#400 gamma=32'd3;row=32'd316;
#400 gamma=32'd4;row=32'd432;
#400 gamma=32'd4;row=32'd392;
#400 gamma=32'd1;row=32'd555;
#400 gamma=32'd3;row=32'd308;
#400 gamma=32'd2;row=32'd295;
#400 gamma=32'd3;row=32'd445;
#400 gamma=32'd3;row=32'd173;
#400 gamma=32'd1;row=32'd81;
#400 gamma=32'd3;row=32'd364;
#400 gamma=32'd5;row=32'd501;
#400 gamma=32'd1;row=32'd276;
#400 gamma=32'd5;row=32'd35;
#400 gamma=32'd2;row=32'd209;
#400 gamma=32'd2;row=32'd67;
#400 gamma=32'd3;row=32'd476;
#400 gamma=32'd2;row=32'd382;
#400 gamma=32'd1;row=32'd69;
#400 gamma=32'd5;row=32'd200;
#400 gamma=32'd5;row=32'd455;
#400 gamma=32'd4;row=32'd438;
#400 gamma=32'd2;row=32'd481;
#400 gamma=32'd4;row=32'd288;
#400 gamma=32'd3;row=32'd521;
#400 gamma=32'd3;row=32'd267;
#400 gamma=32'd2;row=32'd438;
#400 gamma=32'd1;row=32'd513;
#400 gamma=32'd3;row=32'd262;
#400 gamma=32'd5;row=32'd483;
#400 gamma=32'd4;row=32'd142;
#400 gamma=32'd3;row=32'd188;
#400 gamma=32'd5;row=32'd9;
#400 gamma=32'd5;row=32'd362;
#400 gamma=32'd5;row=32'd559;
#400 gamma=32'd2;row=32'd119;
#400 gamma=32'd2;row=32'd135;
#400 gamma=32'd5;row=32'd17;
#400 gamma=32'd1;row=32'd246;
#400 gamma=32'd3;row=32'd507;
#400 gamma=32'd5;row=32'd194;
#400 gamma=32'd2;row=32'd109;
#400 gamma=32'd2;row=32'd153;
#400 gamma=32'd3;row=32'd426;
#400 gamma=32'd2;row=32'd455;
#400 gamma=32'd3;row=32'd429;
#400 gamma=32'd3;row=32'd509;
#400 gamma=32'd1;row=32'd94;
#400 gamma=32'd5;row=32'd387;
#400 gamma=32'd2;row=32'd191;
#400 gamma=32'd2;row=32'd324;
#400 gamma=32'd2;row=32'd266;
#400 gamma=32'd3;row=32'd15;
#400 gamma=32'd4;row=32'd83;
#400 gamma=32'd1;row=32'd19;
#400 gamma=32'd5;row=32'd231;
#400 gamma=32'd3;row=32'd405;
#400 gamma=32'd5;row=32'd543;
#400 gamma=32'd4;row=32'd432;
#400 gamma=32'd1;row=32'd334;
#400 gamma=32'd4;row=32'd456;
#400 gamma=32'd4;row=32'd505;
#400 gamma=32'd5;row=32'd41;
#400 gamma=32'd2;row=32'd123;
#400 gamma=32'd5;row=32'd372;
#400 gamma=32'd1;row=32'd374;
#400 gamma=32'd2;row=32'd152;
#400 gamma=32'd3;row=32'd30;
#400 gamma=32'd4;row=32'd53;
#400 gamma=32'd1;row=32'd189;
#400 gamma=32'd2;row=32'd3;
#400 gamma=32'd5;row=32'd269;
#400 gamma=32'd4;row=32'd221;
#400 gamma=32'd5;row=32'd361;
#400 gamma=32'd5;row=32'd419;
#400 gamma=32'd4;row=32'd112;
#400 gamma=32'd4;row=32'd185;
#400 gamma=32'd3;row=32'd106;
#400 gamma=32'd5;row=32'd351;
#400 gamma=32'd4;row=32'd530;
#400 gamma=32'd2;row=32'd327;
#400 gamma=32'd3;row=32'd40;
#400 gamma=32'd4;row=32'd266;
#400 gamma=32'd1;row=32'd310;
#400 gamma=32'd5;row=32'd19;
#400 gamma=32'd3;row=32'd428;
#400 gamma=32'd3;row=32'd189;
#400 gamma=32'd1;row=32'd479;
#400 gamma=32'd1;row=32'd446;
#400 gamma=32'd5;row=32'd440;
#400 gamma=32'd1;row=32'd96;
#400 gamma=32'd2;row=32'd32;
#400 gamma=32'd5;row=32'd253;
#400 gamma=32'd4;row=32'd242;
#400 gamma=32'd4;row=32'd72;
#400 gamma=32'd1;row=32'd371;
#400 gamma=32'd2;row=32'd265;
#400 gamma=32'd5;row=32'd441;
#400 gamma=32'd3;row=32'd431;
#400 gamma=32'd3;row=32'd524;
#400 gamma=32'd5;row=32'd536;
#400 gamma=32'd2;row=32'd278;
#400 gamma=32'd4;row=32'd334;
#400 gamma=32'd4;row=32'd357;
#400 gamma=32'd3;row=32'd280;
#400 gamma=32'd2;row=32'd285;
#400 gamma=32'd5;row=32'd310;
#400 gamma=32'd2;row=32'd329;
#400 gamma=32'd1;row=32'd415;
#400 gamma=32'd3;row=32'd464;
#400 gamma=32'd3;row=32'd179;
#400 gamma=32'd4;row=32'd53;
#400 gamma=32'd5;row=32'd432;
#400 gamma=32'd5;row=32'd21;
#400 gamma=32'd5;row=32'd476;
#400 gamma=32'd2;row=32'd474;
#400 gamma=32'd1;row=32'd285;
#400 gamma=32'd3;row=32'd202;
#400 gamma=32'd4;row=32'd495;
#400 gamma=32'd4;row=32'd553;
#400 gamma=32'd1;row=32'd544;
#400 gamma=32'd1;row=32'd80;
#400 gamma=32'd4;row=32'd535;
#400 gamma=32'd4;row=32'd288;
#400 gamma=32'd1;row=32'd278;
#400 gamma=32'd1;row=32'd4;
#400 gamma=32'd3;row=32'd28;
#400 gamma=32'd1;row=32'd150;
#400 gamma=32'd2;row=32'd451;
#400 gamma=32'd3;row=32'd349;
#400 gamma=32'd3;row=32'd235;
#400 gamma=32'd1;row=32'd529;
#400 gamma=32'd4;row=32'd99;
#400 gamma=32'd5;row=32'd234;
#400 gamma=32'd3;row=32'd413;
#400 gamma=32'd1;row=32'd250;
#400 gamma=32'd5;row=32'd84;
#400 gamma=32'd4;row=32'd44;
#400 gamma=32'd2;row=32'd505;
#400 gamma=32'd1;row=32'd240;
#400 gamma=32'd2;row=32'd169;
#400 gamma=32'd3;row=32'd388;
#400 gamma=32'd3;row=32'd1;
#400 gamma=32'd5;row=32'd50;
#400 gamma=32'd4;row=32'd93;
#400 gamma=32'd2;row=32'd115;
#400 gamma=32'd5;row=32'd539;
#400 gamma=32'd3;row=32'd296;
#400 gamma=32'd3;row=32'd396;
#400 gamma=32'd5;row=32'd12;
#400 gamma=32'd4;row=32'd10;
#400 gamma=32'd1;row=32'd389;
#400 gamma=32'd4;row=32'd294;
#400 gamma=32'd5;row=32'd470;
#400 gamma=32'd2;row=32'd196;
#400 gamma=32'd3;row=32'd110;
#400 gamma=32'd4;row=32'd202;
#400 gamma=32'd1;row=32'd513;
#400 gamma=32'd2;row=32'd292;
#400 gamma=32'd2;row=32'd289;
#400 gamma=32'd5;row=32'd220;
#400 gamma=32'd2;row=32'd498;
#400 gamma=32'd3;row=32'd316;
#400 gamma=32'd3;row=32'd96;
#400 gamma=32'd5;row=32'd221;
#400 gamma=32'd3;row=32'd214;
#400 gamma=32'd4;row=32'd401;
#400 gamma=32'd1;row=32'd65;
#400 gamma=32'd2;row=32'd220;
#400 gamma=32'd1;row=32'd30;
#400 gamma=32'd5;row=32'd439;
#400 gamma=32'd1;row=32'd41;
#400 gamma=32'd2;row=32'd524;
#400 gamma=32'd2;row=32'd485;
#400 gamma=32'd3;row=32'd300;
#400 gamma=32'd1;row=32'd50;
#400 gamma=32'd5;row=32'd232;
#400 gamma=32'd3;row=32'd205;
#400 gamma=32'd3;row=32'd542;
#400 gamma=32'd2;row=32'd339;
#400 gamma=32'd2;row=32'd188;
#400 gamma=32'd2;row=32'd61;
#400 gamma=32'd2;row=32'd39;
#400 gamma=32'd1;row=32'd511;
#400 gamma=32'd1;row=32'd297;
#400 gamma=32'd2;row=32'd462;
#400 gamma=32'd1;row=32'd144;
#400 gamma=32'd4;row=32'd164;
#400 gamma=32'd2;row=32'd419;
#400 gamma=32'd2;row=32'd253;
#400 gamma=32'd4;row=32'd166;
#400 gamma=32'd4;row=32'd188;
#400 gamma=32'd1;row=32'd478;
#400 gamma=32'd5;row=32'd63;
#400 gamma=32'd3;row=32'd87;
#400 gamma=32'd2;row=32'd320;
#400 gamma=32'd2;row=32'd309;
#400 gamma=32'd2;row=32'd128;
#400 gamma=32'd4;row=32'd203;
#400 gamma=32'd2;row=32'd545;
#400 gamma=32'd1;row=32'd286;
#400 gamma=32'd3;row=32'd296;
#400 gamma=32'd1;row=32'd414;
#400 gamma=32'd5;row=32'd170;
#400 gamma=32'd2;row=32'd538;
#400 gamma=32'd2;row=32'd224;
#400 gamma=32'd1;row=32'd272;
#400 gamma=32'd1;row=32'd362;
#400 gamma=32'd5;row=32'd310;
#400 gamma=32'd3;row=32'd241;
#400 gamma=32'd2;row=32'd133;
#400 gamma=32'd4;row=32'd41;
#400 gamma=32'd2;row=32'd158;
#400 gamma=32'd3;row=32'd488;
#400 gamma=32'd3;row=32'd463;
#400 gamma=32'd5;row=32'd231;
#400 gamma=32'd2;row=32'd364;
#400 gamma=32'd1;row=32'd436;
#400 gamma=32'd5;row=32'd522;
#400 gamma=32'd5;row=32'd372;
#400 gamma=32'd2;row=32'd287;
#400 gamma=32'd1;row=32'd265;
#400 gamma=32'd1;row=32'd555;
#400 gamma=32'd1;row=32'd239;
#400 gamma=32'd3;row=32'd474;
#400 gamma=32'd1;row=32'd371;
#400 gamma=32'd3;row=32'd557;
#400 gamma=32'd2;row=32'd257;
#400 gamma=32'd2;row=32'd361;
#400 gamma=32'd2;row=32'd358;
#400 gamma=32'd3;row=32'd131;
#400 gamma=32'd5;row=32'd259;
#400 gamma=32'd3;row=32'd409;
#400 gamma=32'd4;row=32'd422;
#400 gamma=32'd3;row=32'd111;
#400 gamma=32'd3;row=32'd353;
#400 gamma=32'd2;row=32'd63;
#400 gamma=32'd1;row=32'd531;
#400 gamma=32'd4;row=32'd24;
#400 gamma=32'd5;row=32'd359;
#400 gamma=32'd4;row=32'd414;
#400 gamma=32'd2;row=32'd396;
#400 gamma=32'd1;row=32'd551;
#400 gamma=32'd5;row=32'd167;
#400 gamma=32'd3;row=32'd392;
#400 gamma=32'd5;row=32'd348;
#400 gamma=32'd5;row=32'd78;
#400 gamma=32'd5;row=32'd60;
#400 gamma=32'd5;row=32'd360;
#400 gamma=32'd3;row=32'd53;
#400 gamma=32'd1;row=32'd483;
#400 gamma=32'd4;row=32'd420;
#400 gamma=32'd2;row=32'd246;
#400 gamma=32'd3;row=32'd115;
#400 gamma=32'd2;row=32'd73;
#400 gamma=32'd1;row=32'd152;
#400 gamma=32'd5;row=32'd254;
#400 gamma=32'd2;row=32'd44;
#400 gamma=32'd3;row=32'd383;
#400 gamma=32'd5;row=32'd26;
#400 gamma=32'd2;row=32'd188;
#400 gamma=32'd3;row=32'd427;
#400 gamma=32'd1;row=32'd75;
#400 gamma=32'd3;row=32'd240;
#400 gamma=32'd4;row=32'd423;
#400 gamma=32'd4;row=32'd216;
#400 gamma=32'd3;row=32'd435;
#400 gamma=32'd1;row=32'd246;
#400 gamma=32'd4;row=32'd218;
#400 gamma=32'd5;row=32'd140;
#400 gamma=32'd3;row=32'd109;
#400 gamma=32'd5;row=32'd309;
#400 gamma=32'd3;row=32'd194;
#400 gamma=32'd3;row=32'd315;
#400 gamma=32'd3;row=32'd2;
#400 gamma=32'd3;row=32'd160;
#400 gamma=32'd1;row=32'd189;
#400 gamma=32'd2;row=32'd83;
#400 gamma=32'd5;row=32'd91;
#400 gamma=32'd1;row=32'd153;
#400 gamma=32'd4;row=32'd525;
#400 gamma=32'd5;row=32'd168;
#400 gamma=32'd5;row=32'd27;
#400 gamma=32'd3;row=32'd281;
#400 gamma=32'd3;row=32'd505;
#400 gamma=32'd5;row=32'd225;
#400 gamma=32'd1;row=32'd126;
#400 gamma=32'd5;row=32'd244;
#400 gamma=32'd2;row=32'd323;
#400 gamma=32'd4;row=32'd20;
#400 gamma=32'd5;row=32'd231;
#400 gamma=32'd4;row=32'd4;
#400 gamma=32'd1;row=32'd223;
#400 gamma=32'd4;row=32'd132;
#400 gamma=32'd2;row=32'd182;
#400 gamma=32'd2;row=32'd87;
#400 gamma=32'd4;row=32'd145;
#400 gamma=32'd3;row=32'd461;
#400 gamma=32'd3;row=32'd278;
#400 gamma=32'd5;row=32'd20;
#400 gamma=32'd5;row=32'd341;
#400 gamma=32'd3;row=32'd279;
#400 gamma=32'd4;row=32'd255;
#400 gamma=32'd3;row=32'd488;
#400 gamma=32'd5;row=32'd258;
#400 gamma=32'd1;row=32'd407;
#400 gamma=32'd5;row=32'd289;
#400 gamma=32'd1;row=32'd144;
#400 gamma=32'd2;row=32'd467;
#400 gamma=32'd5;row=32'd154;
#400 gamma=32'd5;row=32'd90;
#400 gamma=32'd3;row=32'd112;
#400 gamma=32'd3;row=32'd466;
#400 gamma=32'd2;row=32'd114;
#400 gamma=32'd2;row=32'd122;
#400 gamma=32'd4;row=32'd415;
#400 gamma=32'd3;row=32'd12;
#400 gamma=32'd2;row=32'd91;
#400 gamma=32'd1;row=32'd114;
#400 gamma=32'd5;row=32'd361;
#400 gamma=32'd1;row=32'd149;
#400 gamma=32'd2;row=32'd25;
#400 gamma=32'd1;row=32'd242;
#400 gamma=32'd2;row=32'd307;
#400 gamma=32'd2;row=32'd485;
#400 gamma=32'd3;row=32'd77;
#400 gamma=32'd1;row=32'd166;
#400 gamma=32'd1;row=32'd404;
#400 gamma=32'd4;row=32'd454;
#400 gamma=32'd4;row=32'd421;
#400 gamma=32'd1;row=32'd495;
#400 gamma=32'd3;row=32'd362;
#400 gamma=32'd2;row=32'd455;
#400 gamma=32'd5;row=32'd17;
#400 gamma=32'd5;row=32'd326;
#400 gamma=32'd1;row=32'd161;
#400 gamma=32'd2;row=32'd387;
#400 gamma=32'd3;row=32'd174;
#400 gamma=32'd5;row=32'd471;
#400 gamma=32'd4;row=32'd337;
#400 gamma=32'd1;row=32'd70;
#400 gamma=32'd1;row=32'd470;
#400 gamma=32'd5;row=32'd246;
#400 gamma=32'd1;row=32'd289;
#400 gamma=32'd1;row=32'd213;
#400 gamma=32'd3;row=32'd480;
#400 gamma=32'd3;row=32'd104;
#400 gamma=32'd1;row=32'd11;
#400 gamma=32'd4;row=32'd172;
#400 gamma=32'd3;row=32'd281;
#400 gamma=32'd4;row=32'd531;
#400 gamma=32'd5;row=32'd220;
#400 gamma=32'd3;row=32'd150;
#400 gamma=32'd1;row=32'd231;
#400 gamma=32'd1;row=32'd381;
#400 gamma=32'd5;row=32'd83;
#400 gamma=32'd3;row=32'd280;
#400 gamma=32'd1;row=32'd528;
#400 gamma=32'd1;row=32'd340;
#400 gamma=32'd2;row=32'd397;
#400 gamma=32'd2;row=32'd294;
#400 gamma=32'd2;row=32'd175;
#400 gamma=32'd3;row=32'd485;
#400 gamma=32'd4;row=32'd340;
#400 gamma=32'd2;row=32'd81;
#400 gamma=32'd1;row=32'd456;
#400 gamma=32'd4;row=32'd550;
#400 gamma=32'd5;row=32'd200;
#400 gamma=32'd5;row=32'd2;
#400 gamma=32'd5;row=32'd293;
#400 gamma=32'd5;row=32'd219;
#400 gamma=32'd1;row=32'd299;
#400 gamma=32'd1;row=32'd78;
#400 gamma=32'd2;row=32'd136;
#400 gamma=32'd5;row=32'd399;
#400 gamma=32'd3;row=32'd162;
#400 gamma=32'd4;row=32'd114;
#400 gamma=32'd5;row=32'd33;
#400 gamma=32'd1;row=32'd365;
#400 gamma=32'd3;row=32'd534;
#400 gamma=32'd4;row=32'd484;
#400 gamma=32'd3;row=32'd557;
#400 gamma=32'd1;row=32'd58;
#400 gamma=32'd2;row=32'd399;
#400 gamma=32'd3;row=32'd363;
#400 gamma=32'd1;row=32'd273;
#400 gamma=32'd2;row=32'd524;
#400 gamma=32'd3;row=32'd82;
#400 gamma=32'd2;row=32'd279;
#400 gamma=32'd2;row=32'd131;
#400 gamma=32'd2;row=32'd145;
#400 gamma=32'd4;row=32'd347;
#400 gamma=32'd2;row=32'd233;
#400 gamma=32'd3;row=32'd25;
#400 gamma=32'd4;row=32'd461;
#400 gamma=32'd4;row=32'd497;
#400 gamma=32'd5;row=32'd37;
#400 gamma=32'd3;row=32'd515;
#400 gamma=32'd4;row=32'd541;
#400 gamma=32'd5;row=32'd240;
#400 gamma=32'd5;row=32'd2;
#400 gamma=32'd1;row=32'd305;
#400 gamma=32'd4;row=32'd267;
#400 gamma=32'd1;row=32'd88;
#400 gamma=32'd1;row=32'd228;
#400 gamma=32'd1;row=32'd121;
#400 gamma=32'd5;row=32'd502;
#400 gamma=32'd3;row=32'd522;
#400 gamma=32'd2;row=32'd131;
#400 gamma=32'd5;row=32'd476;
#400 gamma=32'd1;row=32'd319;
#400 gamma=32'd2;row=32'd250;
#400 gamma=32'd2;row=32'd403;
#400 gamma=32'd4;row=32'd459;
#400 gamma=32'd4;row=32'd293;
#400 gamma=32'd4;row=32'd187;
#400 gamma=32'd2;row=32'd497;
#400 gamma=32'd1;row=32'd399;
#400 gamma=32'd5;row=32'd72;
#400 gamma=32'd3;row=32'd529;
#400 gamma=32'd5;row=32'd293;
#400 gamma=32'd5;row=32'd341;
#400 gamma=32'd5;row=32'd198;
#400 gamma=32'd4;row=32'd538;
#400 gamma=32'd4;row=32'd103;
#400 gamma=32'd2;row=32'd177;
#400 gamma=32'd4;row=32'd222;
#400 gamma=32'd4;row=32'd477;
#400 gamma=32'd1;row=32'd407;
#400 gamma=32'd1;row=32'd534;
#400 gamma=32'd3;row=32'd260;
#400 gamma=32'd2;row=32'd461;
#400 gamma=32'd1;row=32'd176;
#400 gamma=32'd1;row=32'd303;
#400 gamma=32'd3;row=32'd417;
#400 gamma=32'd5;row=32'd442;
#400 gamma=32'd5;row=32'd346;
#400 gamma=32'd4;row=32'd83;
#400 gamma=32'd5;row=32'd430;
#400 gamma=32'd3;row=32'd44;
#400 gamma=32'd5;row=32'd445;
#400 gamma=32'd5;row=32'd499;
#400 gamma=32'd2;row=32'd213;
#400 gamma=32'd1;row=32'd185;
#400 gamma=32'd1;row=32'd354;
#400 gamma=32'd5;row=32'd128;
#400 gamma=32'd1;row=32'd350;
#400 gamma=32'd4;row=32'd460;
#400 gamma=32'd3;row=32'd468;
#400 gamma=32'd4;row=32'd160;
#400 gamma=32'd3;row=32'd347;
#400 gamma=32'd1;row=32'd231;
#400 gamma=32'd2;row=32'd45;
#400 gamma=32'd5;row=32'd352;
#400 gamma=32'd1;row=32'd497;
#400 gamma=32'd1;row=32'd147;
#400 gamma=32'd4;row=32'd473;
#400 gamma=32'd1;row=32'd497;
#400 gamma=32'd2;row=32'd1;
#400 gamma=32'd3;row=32'd509;
#400 gamma=32'd1;row=32'd456;
#400 gamma=32'd2;row=32'd354;
#400 gamma=32'd4;row=32'd204;
#400 gamma=32'd1;row=32'd175;
#400 gamma=32'd2;row=32'd530;
#400 gamma=32'd1;row=32'd211;
#400 gamma=32'd1;row=32'd450;
#400 gamma=32'd2;row=32'd14;
#400 gamma=32'd3;row=32'd542;
#400 gamma=32'd1;row=32'd398;
#400 gamma=32'd1;row=32'd360;
#400 gamma=32'd5;row=32'd379;
#400 gamma=32'd3;row=32'd384;
#400 gamma=32'd2;row=32'd288;
#400 gamma=32'd4;row=32'd436;
#400 gamma=32'd1;row=32'd527;
#400 gamma=32'd4;row=32'd20;
#400 gamma=32'd4;row=32'd102;
#400 gamma=32'd3;row=32'd171;
#400 gamma=32'd1;row=32'd473;
#400 gamma=32'd1;row=32'd396;
#400 gamma=32'd1;row=32'd333;
#400 gamma=32'd3;row=32'd280;
#400 gamma=32'd4;row=32'd22;
#400 gamma=32'd5;row=32'd106;
#400 gamma=32'd1;row=32'd133;
#400 gamma=32'd3;row=32'd501;
#400 gamma=32'd4;row=32'd482;
#400 gamma=32'd2;row=32'd16;
#400 gamma=32'd4;row=32'd485;
#400 gamma=32'd5;row=32'd269;
#400 gamma=32'd5;row=32'd166;
#400 gamma=32'd3;row=32'd88;
#400 gamma=32'd3;row=32'd367;
#400 gamma=32'd1;row=32'd489;
#400 gamma=32'd2;row=32'd175;
#400 gamma=32'd2;row=32'd46;
#400 gamma=32'd1;row=32'd157;
#400 gamma=32'd5;row=32'd358;
#400 gamma=32'd2;row=32'd139;
#400 gamma=32'd3;row=32'd134;
#400 gamma=32'd3;row=32'd434;
#400 gamma=32'd4;row=32'd339;
#400 gamma=32'd3;row=32'd128;
#400 gamma=32'd4;row=32'd355;
#400 gamma=32'd2;row=32'd29;
#400 gamma=32'd5;row=32'd506;
#400 gamma=32'd4;row=32'd191;
#400 gamma=32'd2;row=32'd113;
#400 gamma=32'd3;row=32'd249;
#400 gamma=32'd4;row=32'd523;
#400 gamma=32'd4;row=32'd114;
#400 gamma=32'd1;row=32'd72;
#400 gamma=32'd2;row=32'd358;
#400 gamma=32'd5;row=32'd152;
#400 gamma=32'd5;row=32'd319;
#400 gamma=32'd2;row=32'd209;
#400 gamma=32'd1;row=32'd368;
#400 gamma=32'd2;row=32'd440;
#400 gamma=32'd3;row=32'd19;
#400 gamma=32'd5;row=32'd67;
#400 gamma=32'd2;row=32'd50;
#400 gamma=32'd3;row=32'd497;
#400 gamma=32'd5;row=32'd24;
#400 gamma=32'd1;row=32'd136;
#400 gamma=32'd5;row=32'd121;
#400 gamma=32'd1;row=32'd329;
#400 gamma=32'd1;row=32'd448;
#400 gamma=32'd5;row=32'd223;
#400 gamma=32'd1;row=32'd322;
#400 gamma=32'd2;row=32'd246;
#400 gamma=32'd2;row=32'd136;
#400 gamma=32'd1;row=32'd275;
#400 gamma=32'd3;row=32'd142;
#400 gamma=32'd3;row=32'd505;
#400 gamma=32'd1;row=32'd202;
#400 gamma=32'd3;row=32'd69;
#400 gamma=32'd3;row=32'd207;
#400 gamma=32'd2;row=32'd443;
#400 gamma=32'd2;row=32'd552;
#400 gamma=32'd2;row=32'd403;
#400 gamma=32'd4;row=32'd535;
#400 gamma=32'd5;row=32'd288;
#400 gamma=32'd3;row=32'd180;
#400 gamma=32'd1;row=32'd422;
#400 gamma=32'd5;row=32'd364;
#400 gamma=32'd3;row=32'd527;
#400 gamma=32'd5;row=32'd305;
#400 gamma=32'd5;row=32'd477;
#400 gamma=32'd3;row=32'd23;
#400 gamma=32'd3;row=32'd411;
#400 gamma=32'd2;row=32'd222;
#400 gamma=32'd4;row=32'd12;
#400 gamma=32'd2;row=32'd558;
#400 gamma=32'd1;row=32'd347;
#400 gamma=32'd1;row=32'd385;
#400 gamma=32'd1;row=32'd55;
#400 gamma=32'd3;row=32'd460;
#400 gamma=32'd5;row=32'd181;
#400 gamma=32'd2;row=32'd62;
#400 gamma=32'd4;row=32'd111;
#400 gamma=32'd1;row=32'd81;
#400 gamma=32'd1;row=32'd296;
#400 gamma=32'd1;row=32'd495;
#400 gamma=32'd5;row=32'd517;
#400 gamma=32'd5;row=32'd11;
#400 gamma=32'd4;row=32'd224;
#400 gamma=32'd3;row=32'd237;
#400 gamma=32'd3;row=32'd548;
#400 gamma=32'd2;row=32'd310;
#400 gamma=32'd2;row=32'd28;
#400 gamma=32'd1;row=32'd292;
#400 gamma=32'd4;row=32'd265;
#400 gamma=32'd5;row=32'd419;
#400 gamma=32'd5;row=32'd28;
#400 gamma=32'd3;row=32'd352;
#400 gamma=32'd1;row=32'd133;
#400 gamma=32'd1;row=32'd397;
#400 gamma=32'd2;row=32'd271;
#400 gamma=32'd5;row=32'd308;
#400 gamma=32'd2;row=32'd204;
#400 gamma=32'd4;row=32'd31;
#400 gamma=32'd5;row=32'd50;
#400 gamma=32'd1;row=32'd80;
#400 gamma=32'd5;row=32'd316;
#400 gamma=32'd4;row=32'd110;
#400 gamma=32'd2;row=32'd29;
#400 gamma=32'd3;row=32'd2;
#400 gamma=32'd4;row=32'd201;
#400 gamma=32'd3;row=32'd161;
#400 gamma=32'd5;row=32'd290;
#400 gamma=32'd3;row=32'd300;
#400 gamma=32'd1;row=32'd89;
#400 gamma=32'd5;row=32'd478;
#400 gamma=32'd2;row=32'd521;
#400 gamma=32'd5;row=32'd133;
#400 gamma=32'd2;row=32'd553;
#400 gamma=32'd1;row=32'd477;
#400 gamma=32'd3;row=32'd549;
#400 gamma=32'd5;row=32'd0;
#400 gamma=32'd2;row=32'd189;
#400 gamma=32'd4;row=32'd381;
#400 gamma=32'd3;row=32'd141;
#400 gamma=32'd2;row=32'd471;
#400 gamma=32'd3;row=32'd250;
#400 gamma=32'd1;row=32'd152;
#400 gamma=32'd5;row=32'd252;
#400 gamma=32'd3;row=32'd242;
#400 gamma=32'd2;row=32'd530;
#400 gamma=32'd1;row=32'd165;
#400 gamma=32'd4;row=32'd74;
#400 gamma=32'd4;row=32'd107;
#400 gamma=32'd3;row=32'd390;
#400 gamma=32'd3;row=32'd123;
#400 gamma=32'd5;row=32'd87;
#400 gamma=32'd2;row=32'd545;
#400 gamma=32'd2;row=32'd326;
#400 gamma=32'd2;row=32'd516;
#400 gamma=32'd4;row=32'd232;
#400 gamma=32'd5;row=32'd359;
#400 gamma=32'd5;row=32'd368;
#400 gamma=32'd2;row=32'd342;
#400 gamma=32'd2;row=32'd454;
#400 gamma=32'd2;row=32'd88;
#400 gamma=32'd1;row=32'd38;
#400 gamma=32'd3;row=32'd534;
#400 gamma=32'd5;row=32'd5;
#400 gamma=32'd4;row=32'd458;
#400 gamma=32'd3;row=32'd546;
#400 gamma=32'd4;row=32'd502;
#400 gamma=32'd3;row=32'd372;
#400 gamma=32'd4;row=32'd268;
#400 gamma=32'd4;row=32'd168;
#400 gamma=32'd4;row=32'd495;
#400 gamma=32'd4;row=32'd117;
#400 gamma=32'd1;row=32'd217;
#400 gamma=32'd4;row=32'd204;
#400 gamma=32'd3;row=32'd95;
#400 gamma=32'd1;row=32'd406;
#400 gamma=32'd3;row=32'd393;
#400 gamma=32'd4;row=32'd218;
#400 gamma=32'd2;row=32'd402;
#400 gamma=32'd3;row=32'd243;
#400 gamma=32'd5;row=32'd191;
#400 gamma=32'd2;row=32'd291;
#400 gamma=32'd1;row=32'd132;
#400 gamma=32'd5;row=32'd195;
#400 gamma=32'd5;row=32'd113;
#400 gamma=32'd5;row=32'd512;
#400 gamma=32'd5;row=32'd354;
#400 gamma=32'd5;row=32'd558;
#400 gamma=32'd2;row=32'd425;
#400 gamma=32'd1;row=32'd486;
#400 gamma=32'd5;row=32'd77;
#400 gamma=32'd3;row=32'd439;
#400 gamma=32'd1;row=32'd202;
#400 gamma=32'd1;row=32'd132;
#400 gamma=32'd3;row=32'd366;
#400 gamma=32'd1;row=32'd42;
#400 gamma=32'd1;row=32'd76;
#400 gamma=32'd2;row=32'd367;
#400 gamma=32'd2;row=32'd484;
#400 gamma=32'd2;row=32'd354;
#400 gamma=32'd2;row=32'd503;
#400 gamma=32'd5;row=32'd62;
#400 gamma=32'd2;row=32'd351;
#400 gamma=32'd4;row=32'd481;
#400 gamma=32'd1;row=32'd1;
#400 gamma=32'd1;row=32'd385;
#400 gamma=32'd4;row=32'd432;
#400 gamma=32'd1;row=32'd233;
#400 gamma=32'd5;row=32'd279;
#400 gamma=32'd5;row=32'd361;
#400 gamma=32'd3;row=32'd259;
#400 gamma=32'd4;row=32'd179;
#400 gamma=32'd4;row=32'd555;
#400 gamma=32'd2;row=32'd208;
#400 gamma=32'd2;row=32'd520;
#400 gamma=32'd1;row=32'd558;
#400 gamma=32'd2;row=32'd377;
#400 gamma=32'd3;row=32'd201;
#400 gamma=32'd2;row=32'd316;
#400 gamma=32'd2;row=32'd495;
#400 gamma=32'd3;row=32'd286;
#400 gamma=32'd4;row=32'd502;
#400 gamma=32'd2;row=32'd341;
#400 gamma=32'd3;row=32'd265;
#400 gamma=32'd4;row=32'd237;
#400 gamma=32'd3;row=32'd22;
#400 gamma=32'd2;row=32'd519;
#400 gamma=32'd5;row=32'd110;
#400 gamma=32'd5;row=32'd101;
#400 gamma=32'd3;row=32'd558;
#400 gamma=32'd1;row=32'd414;
#400 gamma=32'd3;row=32'd118;
#400 gamma=32'd4;row=32'd125;
#400 gamma=32'd5;row=32'd88;
#400 gamma=32'd2;row=32'd374;
#400 gamma=32'd3;row=32'd280;
#400 gamma=32'd1;row=32'd136;
#400 gamma=32'd4;row=32'd357;
#400 gamma=32'd2;row=32'd384;
#400 gamma=32'd1;row=32'd391;
#400 gamma=32'd5;row=32'd115;
#400 gamma=32'd4;row=32'd262;
#400 gamma=32'd5;row=32'd129;
#400 gamma=32'd2;row=32'd557;
#400 gamma=32'd2;row=32'd150;
#400 gamma=32'd1;row=32'd397;
#400 gamma=32'd2;row=32'd144;
#400 gamma=32'd1;row=32'd492;
#400 gamma=32'd1;row=32'd446;
#400 gamma=32'd3;row=32'd303;
#400 gamma=32'd3;row=32'd237;
#400 gamma=32'd3;row=32'd333;
#400 gamma=32'd4;row=32'd419;
#400 gamma=32'd1;row=32'd102;
#400 gamma=32'd4;row=32'd423;
#400 gamma=32'd1;row=32'd121;
#400 gamma=32'd5;row=32'd297;
#400 gamma=32'd4;row=32'd515;
#400 gamma=32'd5;row=32'd205;
#400 gamma=32'd4;row=32'd306;
#400 gamma=32'd5;row=32'd34;
#400 gamma=32'd5;row=32'd309;
#400 gamma=32'd2;row=32'd418;
#400 gamma=32'd1;row=32'd396;
#400 gamma=32'd1;row=32'd267;
#400 gamma=32'd4;row=32'd149;
#400 gamma=32'd2;row=32'd318;
#400 gamma=32'd1;row=32'd336;
#400 gamma=32'd1;row=32'd190;
#400 gamma=32'd1;row=32'd43;
#400 gamma=32'd2;row=32'd51;
#400 gamma=32'd3;row=32'd515;
#400 gamma=32'd2;row=32'd106;
#400 gamma=32'd1;row=32'd458;
#400 gamma=32'd1;row=32'd541;
#400 gamma=32'd2;row=32'd464;
#400 gamma=32'd2;row=32'd183;
#400 gamma=32'd5;row=32'd423;
#400 gamma=32'd2;row=32'd273;
#400 gamma=32'd5;row=32'd272;
#400 gamma=32'd1;row=32'd182;
#400 gamma=32'd1;row=32'd479;
#400 gamma=32'd3;row=32'd449;
#400 gamma=32'd3;row=32'd175;
#400 gamma=32'd4;row=32'd361;
#400 gamma=32'd5;row=32'd11;
#400 gamma=32'd1;row=32'd373;
#400 gamma=32'd1;row=32'd479;
#400 gamma=32'd4;row=32'd86;
#400 gamma=32'd3;row=32'd249;
#400 gamma=32'd2;row=32'd352;
#400 gamma=32'd1;row=32'd178;
#400 gamma=32'd1;row=32'd547;
#400 gamma=32'd2;row=32'd354;
#400 gamma=32'd4;row=32'd413;
#400 gamma=32'd3;row=32'd444;
#400 gamma=32'd3;row=32'd72;
#400 gamma=32'd3;row=32'd78;
#400 gamma=32'd2;row=32'd283;
#400 gamma=32'd2;row=32'd105;
#400 gamma=32'd3;row=32'd207;
#400 gamma=32'd3;row=32'd537;
#400 gamma=32'd2;row=32'd237;
#400 gamma=32'd2;row=32'd350;
#400 gamma=32'd4;row=32'd315;
#400 gamma=32'd1;row=32'd414;
#400 gamma=32'd5;row=32'd185;
#400 gamma=32'd2;row=32'd273;
#400 gamma=32'd2;row=32'd164;
#400 gamma=32'd2;row=32'd312;
#400 gamma=32'd4;row=32'd344;
#400 gamma=32'd5;row=32'd275;
#400 gamma=32'd4;row=32'd383;
#400 gamma=32'd2;row=32'd270;
#400 gamma=32'd3;row=32'd244;
#400 gamma=32'd2;row=32'd312;
#400 gamma=32'd2;row=32'd168;
#400 gamma=32'd2;row=32'd542;
#400 gamma=32'd5;row=32'd360;
#400 gamma=32'd3;row=32'd45;
#400 gamma=32'd3;row=32'd299;
#400 gamma=32'd2;row=32'd145;
#400 gamma=32'd1;row=32'd479;
#400 gamma=32'd2;row=32'd47;
#400 gamma=32'd1;row=32'd217;
#400 gamma=32'd3;row=32'd163;
#400 gamma=32'd4;row=32'd3;
#400 gamma=32'd2;row=32'd391;
#400 gamma=32'd4;row=32'd481;
#400 gamma=32'd5;row=32'd67;
#400 gamma=32'd2;row=32'd333;
#400 gamma=32'd2;row=32'd70;
#400 gamma=32'd1;row=32'd55;
#400 gamma=32'd3;row=32'd134;
#400 gamma=32'd5;row=32'd456;
#400 gamma=32'd3;row=32'd304;
#400 gamma=32'd3;row=32'd393;
#400 gamma=32'd4;row=32'd273;
#400 gamma=32'd4;row=32'd90;
#400 gamma=32'd2;row=32'd394;
#400 gamma=32'd3;row=32'd306;
#400 gamma=32'd4;row=32'd110;
#400 gamma=32'd4;row=32'd325;
#400 gamma=32'd1;row=32'd84;
#400 gamma=32'd3;row=32'd51;
#400 gamma=32'd4;row=32'd543;
#400 gamma=32'd3;row=32'd407;
#400 gamma=32'd4;row=32'd76;
#400 gamma=32'd4;row=32'd245;
#400 gamma=32'd4;row=32'd201;
#400 gamma=32'd2;row=32'd515;
#400 gamma=32'd5;row=32'd320;
#400 gamma=32'd5;row=32'd477;
#400 gamma=32'd2;row=32'd28;
#400 gamma=32'd1;row=32'd487;
#400 gamma=32'd5;row=32'd215;
#400 gamma=32'd1;row=32'd396;
#400 gamma=32'd4;row=32'd388;
#400 gamma=32'd5;row=32'd53;
#400 gamma=32'd1;row=32'd173;
#400 gamma=32'd4;row=32'd357;
#400 gamma=32'd3;row=32'd215;
#400 gamma=32'd3;row=32'd555;
#400 gamma=32'd4;row=32'd545;
#400 gamma=32'd3;row=32'd188;
#400 gamma=32'd2;row=32'd306;
#400 gamma=32'd3;row=32'd244;
#400 gamma=32'd2;row=32'd422;
#400 gamma=32'd2;row=32'd146;
#400 gamma=32'd1;row=32'd167;
#400 gamma=32'd4;row=32'd66;
#400 gamma=32'd2;row=32'd251;
#400 gamma=32'd2;row=32'd278;
#400 gamma=32'd2;row=32'd450;
#400 gamma=32'd4;row=32'd126;
#400 gamma=32'd3;row=32'd343;
#400 gamma=32'd5;row=32'd407;
#400 gamma=32'd3;row=32'd413;
#400 gamma=32'd2;row=32'd376;
#400 gamma=32'd3;row=32'd383;
#400 gamma=32'd5;row=32'd38;
#400 gamma=32'd3;row=32'd396;
#400 gamma=32'd1;row=32'd484;
#400 gamma=32'd4;row=32'd253;
#400 gamma=32'd5;row=32'd363;
#400 gamma=32'd1;row=32'd382;
#400 gamma=32'd2;row=32'd255;
#400 gamma=32'd4;row=32'd1;
#400 gamma=32'd4;row=32'd198;
#400 gamma=32'd5;row=32'd57;
#400 gamma=32'd2;row=32'd337;
#400 gamma=32'd5;row=32'd217;
#400 gamma=32'd4;row=32'd80;
#400 gamma=32'd2;row=32'd289;
#400 gamma=32'd5;row=32'd388;
#400 gamma=32'd5;row=32'd491;
#400 gamma=32'd4;row=32'd116;
#400 gamma=32'd4;row=32'd418;
#400 gamma=32'd1;row=32'd539;
#400 gamma=32'd5;row=32'd110;
#400 gamma=32'd2;row=32'd107;
#400 gamma=32'd2;row=32'd85;
#400 gamma=32'd1;row=32'd57;
#400 gamma=32'd3;row=32'd295;
#400 gamma=32'd1;row=32'd221;
#400 gamma=32'd4;row=32'd139;
#400 gamma=32'd3;row=32'd91;
#400 gamma=32'd2;row=32'd436;
#400 gamma=32'd2;row=32'd547;
#400 gamma=32'd3;row=32'd427;
#400 gamma=32'd3;row=32'd536;
#400 gamma=32'd5;row=32'd338;
#400 gamma=32'd5;row=32'd223;
#400 gamma=32'd4;row=32'd486;
#400 gamma=32'd4;row=32'd134;
#400 gamma=32'd3;row=32'd84;
#400 gamma=32'd4;row=32'd417;
#400 gamma=32'd4;row=32'd553;
#400 gamma=32'd1;row=32'd1;
#400 gamma=32'd1;row=32'd408;
#400 gamma=32'd1;row=32'd42;
#400 gamma=32'd5;row=32'd296;
#400 gamma=32'd1;row=32'd22;
#400 gamma=32'd5;row=32'd11;
#400 gamma=32'd4;row=32'd373;
#400 gamma=32'd3;row=32'd133;
#400 gamma=32'd1;row=32'd382;
#400 gamma=32'd1;row=32'd101;
#400 gamma=32'd5;row=32'd478;
#400 gamma=32'd2;row=32'd415;
#400 gamma=32'd2;row=32'd46;
#400 gamma=32'd5;row=32'd395;
#400 gamma=32'd3;row=32'd385;
#400 gamma=32'd5;row=32'd498;
#400 gamma=32'd2;row=32'd138;
#400 gamma=32'd5;row=32'd3;
#400 gamma=32'd1;row=32'd360;
#400 gamma=32'd3;row=32'd56;
#400 gamma=32'd5;row=32'd299;
#400 gamma=32'd1;row=32'd252;
#400 gamma=32'd2;row=32'd143;
#400 gamma=32'd1;row=32'd319;
#400 gamma=32'd4;row=32'd6;
#400 gamma=32'd4;row=32'd61;
#400 gamma=32'd1;row=32'd288;
#400 gamma=32'd4;row=32'd249;
#400 gamma=32'd1;row=32'd450;
#400 gamma=32'd3;row=32'd5;
#400 gamma=32'd1;row=32'd241;
#400 gamma=32'd5;row=32'd490;
#400 gamma=32'd2;row=32'd238;
#400 gamma=32'd5;row=32'd447;
#400 gamma=32'd5;row=32'd216;
#400 gamma=32'd5;row=32'd421;
#400 gamma=32'd2;row=32'd261;
#400 gamma=32'd5;row=32'd123;
#400 gamma=32'd3;row=32'd331;
#400 gamma=32'd3;row=32'd384;
#400 gamma=32'd3;row=32'd130;
#400 gamma=32'd4;row=32'd548;
#400 gamma=32'd1;row=32'd83;
#400 gamma=32'd2;row=32'd421;
#400 gamma=32'd1;row=32'd514;
#400 gamma=32'd5;row=32'd202;
#400 gamma=32'd4;row=32'd272;
#400 gamma=32'd4;row=32'd470;
#400 gamma=32'd2;row=32'd102;
#400 gamma=32'd4;row=32'd223;
#400 gamma=32'd4;row=32'd337;
#400 gamma=32'd3;row=32'd50;
#400 gamma=32'd2;row=32'd66;
#400 gamma=32'd3;row=32'd55;
#400 gamma=32'd3;row=32'd389;
#400 gamma=32'd3;row=32'd139;
#400 gamma=32'd3;row=32'd279;
#400 gamma=32'd2;row=32'd103;
#400 gamma=32'd4;row=32'd456;
#400 gamma=32'd2;row=32'd130;
#400 gamma=32'd5;row=32'd41;
#400 gamma=32'd3;row=32'd219;
#400 gamma=32'd1;row=32'd20;
#400 gamma=32'd4;row=32'd354;
#400 gamma=32'd4;row=32'd546;
#400 gamma=32'd1;row=32'd278;
#400 gamma=32'd4;row=32'd286;
#400 gamma=32'd3;row=32'd26;
#400 gamma=32'd4;row=32'd368;
#400 gamma=32'd5;row=32'd118;
#400 gamma=32'd2;row=32'd487;
#400 gamma=32'd4;row=32'd56;
#400 gamma=32'd2;row=32'd432;
#400 gamma=32'd2;row=32'd301;
#400 gamma=32'd5;row=32'd45;
#400 gamma=32'd4;row=32'd434;
#400 gamma=32'd5;row=32'd321;
#400 gamma=32'd1;row=32'd230;
#400 gamma=32'd3;row=32'd458;
#400 gamma=32'd2;row=32'd212;
#400 gamma=32'd5;row=32'd7;
#400 gamma=32'd1;row=32'd411;
#400 gamma=32'd2;row=32'd97;
#400 gamma=32'd1;row=32'd364;
#400 gamma=32'd3;row=32'd316;
#400 gamma=32'd2;row=32'd454;
#400 gamma=32'd2;row=32'd231;
#400 gamma=32'd4;row=32'd286;
#400 gamma=32'd5;row=32'd276;
#400 gamma=32'd4;row=32'd270;
#400 gamma=32'd2;row=32'd246;
#400 gamma=32'd4;row=32'd319;
#400 gamma=32'd3;row=32'd552;
#400 gamma=32'd4;row=32'd413;
#400 gamma=32'd4;row=32'd60;
#400 gamma=32'd2;row=32'd319;
#400 gamma=32'd4;row=32'd159;
#400 gamma=32'd2;row=32'd33;
#400 gamma=32'd4;row=32'd272;
#400 gamma=32'd3;row=32'd112;
#400 gamma=32'd4;row=32'd158;
#400 gamma=32'd3;row=32'd541;
#400 gamma=32'd4;row=32'd332;
#400 gamma=32'd3;row=32'd515;
#400 gamma=32'd2;row=32'd491;
#400 gamma=32'd3;row=32'd95;
#400 gamma=32'd3;row=32'd107;
#400 gamma=32'd2;row=32'd505;
#400 gamma=32'd1;row=32'd22;
#400 gamma=32'd4;row=32'd252;
#400 gamma=32'd3;row=32'd440;
#400 gamma=32'd4;row=32'd111;
#400 gamma=32'd2;row=32'd286;
#400 gamma=32'd5;row=32'd533;
#400 gamma=32'd2;row=32'd292;
#400 gamma=32'd3;row=32'd543;
#400 gamma=32'd1;row=32'd282;
#400 gamma=32'd4;row=32'd137;
#400 gamma=32'd3;row=32'd237;
#400 gamma=32'd4;row=32'd244;
#400 gamma=32'd5;row=32'd256;
#400 gamma=32'd1;row=32'd146;
#400 gamma=32'd2;row=32'd270;
#400 gamma=32'd5;row=32'd299;
#400 gamma=32'd4;row=32'd142;
#400 gamma=32'd5;row=32'd76;
#400 gamma=32'd4;row=32'd124;
#400 gamma=32'd5;row=32'd147;
#400 gamma=32'd4;row=32'd201;
#400 gamma=32'd2;row=32'd497;
#400 gamma=32'd2;row=32'd37;
#400 gamma=32'd4;row=32'd474;
#400 gamma=32'd5;row=32'd413;
#400 gamma=32'd2;row=32'd157;
#400 gamma=32'd3;row=32'd404;
#400 gamma=32'd3;row=32'd202;
#400 gamma=32'd2;row=32'd493;
#400 gamma=32'd5;row=32'd396;
#400 gamma=32'd3;row=32'd523;
#400 gamma=32'd3;row=32'd471;
#400 gamma=32'd2;row=32'd329;
#400 gamma=32'd2;row=32'd553;
#400 gamma=32'd5;row=32'd484;
#400 gamma=32'd2;row=32'd104;
#400 gamma=32'd3;row=32'd204;
#400 gamma=32'd2;row=32'd129;
#400 gamma=32'd5;row=32'd110;
#400 gamma=32'd1;row=32'd286;
#400 gamma=32'd4;row=32'd495;
#400 gamma=32'd4;row=32'd37;
#400 gamma=32'd3;row=32'd0;
#400 gamma=32'd2;row=32'd302;
#400 gamma=32'd5;row=32'd340;
#400 gamma=32'd2;row=32'd418;
#400 gamma=32'd1;row=32'd110;
#400 gamma=32'd1;row=32'd514;
#400 gamma=32'd5;row=32'd485;
#400 gamma=32'd4;row=32'd279;
#400 gamma=32'd4;row=32'd297;
#400 gamma=32'd2;row=32'd176;
#400 gamma=32'd1;row=32'd10;
#400 gamma=32'd2;row=32'd136;
#400 gamma=32'd2;row=32'd410;
#400 gamma=32'd2;row=32'd3;
#400 gamma=32'd4;row=32'd444;
#400 gamma=32'd1;row=32'd496;
#400 gamma=32'd1;row=32'd516;
#400 gamma=32'd4;row=32'd291;
#400 gamma=32'd5;row=32'd203;
#400 gamma=32'd4;row=32'd140;
#400 gamma=32'd3;row=32'd356;
#400 gamma=32'd4;row=32'd55;
#400 gamma=32'd2;row=32'd465;
#400 gamma=32'd1;row=32'd188;
#400 gamma=32'd2;row=32'd547;
#400 gamma=32'd1;row=32'd52;
#400 gamma=32'd3;row=32'd313;
#400 gamma=32'd1;row=32'd98;
#400 gamma=32'd2;row=32'd347;
#400 gamma=32'd1;row=32'd157;
#400 gamma=32'd3;row=32'd159;
#400 gamma=32'd5;row=32'd202;
#400 gamma=32'd5;row=32'd494;
#400 gamma=32'd4;row=32'd194;
#400 gamma=32'd4;row=32'd56;
#400 gamma=32'd1;row=32'd318;
#400 gamma=32'd4;row=32'd510;
#400 gamma=32'd3;row=32'd224;
#400 gamma=32'd1;row=32'd432;
#400 gamma=32'd3;row=32'd556;
#400 gamma=32'd5;row=32'd233;
#400 gamma=32'd2;row=32'd240;
#400 gamma=32'd2;row=32'd139;
#400 gamma=32'd1;row=32'd58;
#400 gamma=32'd5;row=32'd462;
#400 gamma=32'd4;row=32'd406;
#400 gamma=32'd1;row=32'd328;
#400 gamma=32'd4;row=32'd173;
#400 gamma=32'd4;row=32'd141;
#400 gamma=32'd5;row=32'd342;
#400 gamma=32'd3;row=32'd365;
#400 gamma=32'd4;row=32'd360;
#400 gamma=32'd5;row=32'd11;
#400 gamma=32'd4;row=32'd439;
#400 gamma=32'd2;row=32'd127;
#400 gamma=32'd1;row=32'd115;
#400 gamma=32'd3;row=32'd343;
#400 gamma=32'd3;row=32'd456;
#400 gamma=32'd3;row=32'd449;
#400 gamma=32'd3;row=32'd48;
#400 gamma=32'd5;row=32'd283;
#400 gamma=32'd2;row=32'd434;
#400 gamma=32'd2;row=32'd532;
#400 gamma=32'd4;row=32'd19;
#400 gamma=32'd4;row=32'd382;
#400 gamma=32'd4;row=32'd248;
#400 gamma=32'd2;row=32'd82;
#400 gamma=32'd4;row=32'd205;
#400 gamma=32'd2;row=32'd283;
#400 gamma=32'd4;row=32'd102;
#400 gamma=32'd5;row=32'd85;
#400 gamma=32'd3;row=32'd286;
#400 gamma=32'd3;row=32'd523;
#400 gamma=32'd3;row=32'd489;
#400 gamma=32'd5;row=32'd238;
#400 gamma=32'd2;row=32'd315;
#400 gamma=32'd5;row=32'd304;
#400 gamma=32'd2;row=32'd78;
#400 gamma=32'd5;row=32'd246;
#400 gamma=32'd1;row=32'd458;
#400 gamma=32'd2;row=32'd394;
#400 gamma=32'd3;row=32'd366;
#400 gamma=32'd5;row=32'd421;
#400 gamma=32'd3;row=32'd26;
#400 gamma=32'd1;row=32'd417;
#400 gamma=32'd3;row=32'd150;
#400 gamma=32'd2;row=32'd173;
#400 gamma=32'd1;row=32'd517;
#400 gamma=32'd2;row=32'd149;
#400 gamma=32'd3;row=32'd32;
#400 gamma=32'd4;row=32'd71;
#400 gamma=32'd1;row=32'd545;
#400 gamma=32'd5;row=32'd118;
#400 gamma=32'd5;row=32'd179;
#400 gamma=32'd2;row=32'd439;
#400 gamma=32'd5;row=32'd180;
#400 gamma=32'd4;row=32'd188;
#400 gamma=32'd5;row=32'd458;
#400 gamma=32'd4;row=32'd139;
#400 gamma=32'd5;row=32'd441;
#400 gamma=32'd1;row=32'd101;
#400 gamma=32'd4;row=32'd261;
#400 gamma=32'd4;row=32'd204;
#400 gamma=32'd3;row=32'd497;
#400 gamma=32'd5;row=32'd351;
#400 gamma=32'd5;row=32'd391;
#400 gamma=32'd2;row=32'd111;
#400 gamma=32'd5;row=32'd466;
#400 gamma=32'd4;row=32'd193;
#400 gamma=32'd1;row=32'd391;
#400 gamma=32'd4;row=32'd276;
#400 gamma=32'd4;row=32'd536;
#400 gamma=32'd3;row=32'd11;
#400 gamma=32'd1;row=32'd307;
#400 gamma=32'd5;row=32'd263;
#400 gamma=32'd5;row=32'd227;
#400 gamma=32'd1;row=32'd314;
#400 gamma=32'd3;row=32'd48;
#400 gamma=32'd1;row=32'd193;
#400 gamma=32'd3;row=32'd554;
#400 gamma=32'd2;row=32'd558;
#400 gamma=32'd2;row=32'd295;
#400 gamma=32'd4;row=32'd209;
#400 gamma=32'd4;row=32'd353;
#400 gamma=32'd1;row=32'd484;
#400 gamma=32'd2;row=32'd538;
#400 gamma=32'd3;row=32'd436;
#400 gamma=32'd3;row=32'd108;
#400 gamma=32'd3;row=32'd357;
#400 gamma=32'd5;row=32'd72;
#400 gamma=32'd1;row=32'd552;
#400 gamma=32'd2;row=32'd485;
#400 gamma=32'd1;row=32'd150;
#400 gamma=32'd2;row=32'd140;
#400 gamma=32'd4;row=32'd6;
#400 gamma=32'd3;row=32'd250;
#400 gamma=32'd5;row=32'd167;
#400 gamma=32'd5;row=32'd532;
#400 gamma=32'd3;row=32'd341;
#400 gamma=32'd3;row=32'd151;
#400 gamma=32'd2;row=32'd125;
#400 gamma=32'd5;row=32'd431;
#400 gamma=32'd2;row=32'd230;
#400 gamma=32'd3;row=32'd383;
#400 gamma=32'd5;row=32'd442;
#400 gamma=32'd2;row=32'd509;
#400 gamma=32'd2;row=32'd3;
#400 gamma=32'd2;row=32'd211;
#400 gamma=32'd2;row=32'd153;
#400 gamma=32'd5;row=32'd227;
#400 gamma=32'd2;row=32'd260;
#400 gamma=32'd3;row=32'd459;
#400 gamma=32'd3;row=32'd248;
#400 gamma=32'd3;row=32'd43;
#400 gamma=32'd2;row=32'd447;
#400 gamma=32'd1;row=32'd90;
#400 gamma=32'd1;row=32'd148;
#400 gamma=32'd2;row=32'd67;
#400 gamma=32'd4;row=32'd463;
#400 gamma=32'd4;row=32'd295;
#400 gamma=32'd5;row=32'd86;
#400 gamma=32'd2;row=32'd505;
#400 gamma=32'd5;row=32'd516;
#400 gamma=32'd5;row=32'd209;
#400 gamma=32'd2;row=32'd238;
#400 gamma=32'd1;row=32'd374;
#400 gamma=32'd5;row=32'd73;
#400 gamma=32'd5;row=32'd57;
#400 gamma=32'd4;row=32'd537;
#400 gamma=32'd4;row=32'd243;
#400 gamma=32'd5;row=32'd338;
#400 gamma=32'd3;row=32'd31;
#400 gamma=32'd3;row=32'd491;
#400 gamma=32'd3;row=32'd232;
#400 gamma=32'd1;row=32'd353;
#400 gamma=32'd1;row=32'd40;
#400 gamma=32'd4;row=32'd491;
#400 gamma=32'd3;row=32'd182;
#400 gamma=32'd2;row=32'd109;
#400 gamma=32'd2;row=32'd77;
#400 gamma=32'd5;row=32'd292;
#400 gamma=32'd2;row=32'd438;
#400 gamma=32'd4;row=32'd531;
#400 gamma=32'd1;row=32'd236;
#400 gamma=32'd4;row=32'd283;
#400 gamma=32'd2;row=32'd250;
#400 gamma=32'd2;row=32'd281;
#400 gamma=32'd3;row=32'd492;
#400 gamma=32'd5;row=32'd514;
#400 gamma=32'd5;row=32'd167;
#400 gamma=32'd3;row=32'd475;
#400 gamma=32'd4;row=32'd302;
#400 gamma=32'd2;row=32'd100;
#400 gamma=32'd3;row=32'd293;
#400 gamma=32'd2;row=32'd484;
#400 gamma=32'd4;row=32'd196;
#400 gamma=32'd1;row=32'd391;
#400 gamma=32'd2;row=32'd130;
#400 gamma=32'd2;row=32'd21;
#400 gamma=32'd3;row=32'd112;
#400 gamma=32'd1;row=32'd525;
#400 gamma=32'd1;row=32'd552;
#400 gamma=32'd2;row=32'd544;
#400 gamma=32'd1;row=32'd123;
#400 gamma=32'd4;row=32'd423;
#400 gamma=32'd5;row=32'd280;
#400 gamma=32'd5;row=32'd45;
#400 gamma=32'd3;row=32'd95;
#400 gamma=32'd1;row=32'd31;
#400 gamma=32'd3;row=32'd219;
#400 gamma=32'd1;row=32'd108;
#400 gamma=32'd2;row=32'd446;
#400 gamma=32'd5;row=32'd434;
#400 gamma=32'd1;row=32'd147;
#400 gamma=32'd3;row=32'd553;
#400 gamma=32'd5;row=32'd382;
#400 gamma=32'd1;row=32'd136;
#400 gamma=32'd2;row=32'd63;
#400 gamma=32'd5;row=32'd81;
#400 gamma=32'd5;row=32'd126;
#400 gamma=32'd5;row=32'd24;
#400 gamma=32'd1;row=32'd182;
#400 gamma=32'd5;row=32'd64;
#400 gamma=32'd2;row=32'd118;
#400 gamma=32'd2;row=32'd249;
#400 gamma=32'd4;row=32'd394;
#400 gamma=32'd2;row=32'd505;
#400 gamma=32'd1;row=32'd350;
#400 gamma=32'd4;row=32'd444;
#400 gamma=32'd2;row=32'd14;
#400 gamma=32'd5;row=32'd215;
#400 gamma=32'd3;row=32'd419;
#400 gamma=32'd1;row=32'd381;
#400 gamma=32'd2;row=32'd542;
#400 gamma=32'd5;row=32'd222;
#400 gamma=32'd4;row=32'd86;
#400 gamma=32'd5;row=32'd84;
#400 gamma=32'd3;row=32'd435;
#400 gamma=32'd2;row=32'd421;
#400 gamma=32'd1;row=32'd358;
#400 gamma=32'd1;row=32'd495;
#400 gamma=32'd4;row=32'd415;
#400 gamma=32'd4;row=32'd253;
#400 gamma=32'd4;row=32'd458;
#400 gamma=32'd1;row=32'd482;
#400 gamma=32'd3;row=32'd336;
#400 gamma=32'd5;row=32'd26;
#400 gamma=32'd4;row=32'd253;
#400 gamma=32'd4;row=32'd125;
#400 gamma=32'd4;row=32'd4;
#400 gamma=32'd2;row=32'd418;
#400 gamma=32'd3;row=32'd122;
#400 gamma=32'd3;row=32'd257;
#400 gamma=32'd3;row=32'd326;
#400 gamma=32'd2;row=32'd391;
#400 gamma=32'd1;row=32'd293;
#400 gamma=32'd3;row=32'd452;
#400 gamma=32'd4;row=32'd351;
#400 gamma=32'd5;row=32'd33;
#400 gamma=32'd3;row=32'd83;
#400 gamma=32'd5;row=32'd120;
#400 gamma=32'd3;row=32'd558;
#400 gamma=32'd4;row=32'd305;
#400 gamma=32'd2;row=32'd133;
#400 gamma=32'd5;row=32'd201;
#400 gamma=32'd3;row=32'd213;
#400 gamma=32'd4;row=32'd109;
#400 gamma=32'd4;row=32'd445;
#400 gamma=32'd2;row=32'd167;
#400 gamma=32'd1;row=32'd119;
#400 gamma=32'd3;row=32'd359;
#400 gamma=32'd2;row=32'd437;
#400 gamma=32'd5;row=32'd339;
#400 gamma=32'd1;row=32'd537;
#400 gamma=32'd2;row=32'd441;
#400 gamma=32'd5;row=32'd448;
#400 gamma=32'd4;row=32'd529;
#400 gamma=32'd4;row=32'd218;
#400 gamma=32'd3;row=32'd125;
#400 gamma=32'd3;row=32'd338;
#400 gamma=32'd3;row=32'd216;
#400 gamma=32'd5;row=32'd302;
#400 gamma=32'd5;row=32'd180;
#400 gamma=32'd3;row=32'd461;
#400 gamma=32'd5;row=32'd551;
#400 gamma=32'd1;row=32'd498;
#400 gamma=32'd3;row=32'd354;
#400 gamma=32'd5;row=32'd221;
#400 gamma=32'd2;row=32'd51;
#400 gamma=32'd1;row=32'd445;
#400 gamma=32'd5;row=32'd234;
#400 gamma=32'd3;row=32'd425;
#400 gamma=32'd2;row=32'd521;
#400 gamma=32'd1;row=32'd159;
#400 gamma=32'd5;row=32'd285;
#400 gamma=32'd5;row=32'd374;
#400 gamma=32'd5;row=32'd241;
#400 gamma=32'd2;row=32'd379;
#400 gamma=32'd4;row=32'd9;
#400 gamma=32'd3;row=32'd473;
#400 gamma=32'd1;row=32'd538;
#400 gamma=32'd1;row=32'd64;
#400 gamma=32'd5;row=32'd64;
#400 gamma=32'd3;row=32'd319;
#400 gamma=32'd2;row=32'd140;
#400 gamma=32'd4;row=32'd133;
#400 gamma=32'd1;row=32'd108;
#400 gamma=32'd3;row=32'd371;
#400 gamma=32'd3;row=32'd279;
#400 gamma=32'd5;row=32'd8;
#400 gamma=32'd3;row=32'd363;
#400 gamma=32'd3;row=32'd409;
#400 gamma=32'd4;row=32'd328;
#400 gamma=32'd1;row=32'd536;
#400 gamma=32'd4;row=32'd547;
#400 gamma=32'd3;row=32'd444;
#400 gamma=32'd3;row=32'd332;
#400 gamma=32'd5;row=32'd166;
#400 gamma=32'd5;row=32'd253;
#400 gamma=32'd5;row=32'd468;
#400 gamma=32'd3;row=32'd496;
#400 gamma=32'd4;row=32'd124;
#400 gamma=32'd4;row=32'd302;
#400 gamma=32'd3;row=32'd266;
#400 gamma=32'd4;row=32'd403;
#400 gamma=32'd1;row=32'd367;
#400 gamma=32'd1;row=32'd78;
#400 gamma=32'd3;row=32'd296;
#400 gamma=32'd3;row=32'd240;
#400 gamma=32'd1;row=32'd152;
#400 gamma=32'd4;row=32'd387;
#400 gamma=32'd2;row=32'd398;
#400 gamma=32'd1;row=32'd70;
#400 gamma=32'd4;row=32'd452;
#400 gamma=32'd5;row=32'd141;
#400 gamma=32'd2;row=32'd131;
#400 gamma=32'd3;row=32'd460;
#400 gamma=32'd2;row=32'd437;
#400 gamma=32'd5;row=32'd468;
#400 gamma=32'd5;row=32'd76;
#400 gamma=32'd3;row=32'd497;
#400 gamma=32'd3;row=32'd12;
#400 gamma=32'd2;row=32'd534;
#400 gamma=32'd3;row=32'd399;
#400 gamma=32'd2;row=32'd128;
#400 gamma=32'd2;row=32'd50;
#400 gamma=32'd2;row=32'd368;
#400 gamma=32'd5;row=32'd104;
#400 gamma=32'd2;row=32'd365;
#400 gamma=32'd5;row=32'd220;
#400 gamma=32'd4;row=32'd267;
#400 gamma=32'd1;row=32'd156;
#400 gamma=32'd1;row=32'd311;
#400 gamma=32'd5;row=32'd462;
#400 gamma=32'd3;row=32'd255;
#400 gamma=32'd4;row=32'd529;
#400 gamma=32'd5;row=32'd350;
#400 gamma=32'd1;row=32'd4;
#400 gamma=32'd5;row=32'd493;
#400 gamma=32'd1;row=32'd202;
#400 gamma=32'd1;row=32'd529;
#400 gamma=32'd5;row=32'd93;
#400 gamma=32'd1;row=32'd452;
#400 gamma=32'd4;row=32'd532;
#400 gamma=32'd2;row=32'd317;
#400 gamma=32'd4;row=32'd467;
#400 gamma=32'd5;row=32'd424;
#400 gamma=32'd5;row=32'd257;
#400 gamma=32'd3;row=32'd60;
#400 gamma=32'd4;row=32'd428;
#400 gamma=32'd5;row=32'd425;
#400 gamma=32'd3;row=32'd216;
#400 gamma=32'd3;row=32'd294;
#400 gamma=32'd5;row=32'd331;
#400 gamma=32'd5;row=32'd462;
#400 gamma=32'd5;row=32'd494;
#400 gamma=32'd3;row=32'd528;
#400 gamma=32'd1;row=32'd117;
#400 gamma=32'd4;row=32'd399;
#400 gamma=32'd2;row=32'd408;
#400 gamma=32'd4;row=32'd122;
#400 gamma=32'd1;row=32'd27;
#400 gamma=32'd5;row=32'd38;
#400 gamma=32'd2;row=32'd385;
#400 gamma=32'd5;row=32'd65;
#400 gamma=32'd5;row=32'd388;
#400 gamma=32'd1;row=32'd270;
#400 gamma=32'd5;row=32'd263;
#400 gamma=32'd2;row=32'd118;
#400 gamma=32'd2;row=32'd258;
#400 gamma=32'd3;row=32'd11;
#400 gamma=32'd4;row=32'd48;
#400 gamma=32'd4;row=32'd211;
#400 gamma=32'd5;row=32'd445;
#400 gamma=32'd5;row=32'd359;
#400 gamma=32'd1;row=32'd21;
#400 gamma=32'd3;row=32'd47;
#400 gamma=32'd1;row=32'd323;
#400 gamma=32'd4;row=32'd197;
#400 gamma=32'd4;row=32'd359;
#400 gamma=32'd2;row=32'd481;
#400 gamma=32'd4;row=32'd183;
#400 gamma=32'd5;row=32'd354;
#400 gamma=32'd5;row=32'd330;
#400 gamma=32'd3;row=32'd257;
#400 gamma=32'd4;row=32'd358;
#400 gamma=32'd5;row=32'd96;
#400 gamma=32'd1;row=32'd247;
#400 gamma=32'd2;row=32'd182;
#400 gamma=32'd4;row=32'd84;
#400 gamma=32'd4;row=32'd78;
#400 gamma=32'd5;row=32'd139;
#400 gamma=32'd5;row=32'd3;
#400 gamma=32'd2;row=32'd277;
#400 gamma=32'd4;row=32'd147;
#400 gamma=32'd2;row=32'd447;
#400 gamma=32'd3;row=32'd127;
#400 gamma=32'd2;row=32'd0;
#400 gamma=32'd3;row=32'd461;
#400 gamma=32'd3;row=32'd178;
#400 gamma=32'd4;row=32'd428;
#400 gamma=32'd2;row=32'd46;
#400 gamma=32'd4;row=32'd172;
#400 gamma=32'd1;row=32'd364;
#400 gamma=32'd2;row=32'd207;
#400 gamma=32'd2;row=32'd394;
#400 gamma=32'd4;row=32'd266;
#400 gamma=32'd4;row=32'd96;
#400 gamma=32'd1;row=32'd11;
#400 gamma=32'd3;row=32'd48;
#400 gamma=32'd5;row=32'd12;
#400 gamma=32'd5;row=32'd363;
#400 gamma=32'd5;row=32'd477;
#400 gamma=32'd2;row=32'd134;
#400 gamma=32'd3;row=32'd136;
#400 gamma=32'd2;row=32'd113;
#400 gamma=32'd1;row=32'd37;
#400 gamma=32'd4;row=32'd186;
#400 gamma=32'd1;row=32'd214;
#400 gamma=32'd1;row=32'd410;
#400 gamma=32'd2;row=32'd146;
#400 gamma=32'd4;row=32'd473;
#400 gamma=32'd4;row=32'd538;
#400 gamma=32'd2;row=32'd128;
#400 gamma=32'd3;row=32'd187;
#400 gamma=32'd2;row=32'd219;
#400 gamma=32'd5;row=32'd552;
#400 gamma=32'd5;row=32'd311;
#400 gamma=32'd1;row=32'd169;
#400 gamma=32'd5;row=32'd333;
#400 gamma=32'd3;row=32'd88;
#400 gamma=32'd3;row=32'd442;
#400 gamma=32'd1;row=32'd4;
#400 gamma=32'd2;row=32'd498;
#400 gamma=32'd3;row=32'd152;
#400 gamma=32'd3;row=32'd148;
#400 gamma=32'd3;row=32'd222;
#400 gamma=32'd1;row=32'd56;
#400 gamma=32'd4;row=32'd108;
#400 gamma=32'd1;row=32'd524;
#400 gamma=32'd5;row=32'd86;
#400 gamma=32'd3;row=32'd422;
#400 gamma=32'd3;row=32'd176;
#400 gamma=32'd4;row=32'd381;
#400 gamma=32'd3;row=32'd162;
#400 gamma=32'd1;row=32'd352;
#400 gamma=32'd3;row=32'd150;
#400 gamma=32'd3;row=32'd517;
#400 gamma=32'd1;row=32'd264;
#400 gamma=32'd2;row=32'd514;
#400 gamma=32'd3;row=32'd493;
#400 gamma=32'd4;row=32'd299;
#400 gamma=32'd2;row=32'd494;
#400 gamma=32'd2;row=32'd443;
#400 gamma=32'd4;row=32'd320;
#400 gamma=32'd3;row=32'd52;
#400 gamma=32'd3;row=32'd315;
#400 gamma=32'd2;row=32'd456;
#400 gamma=32'd3;row=32'd43;
#400 gamma=32'd2;row=32'd282;
#400 gamma=32'd4;row=32'd152;
#400 gamma=32'd4;row=32'd359;
#400 gamma=32'd1;row=32'd271;
#400 gamma=32'd2;row=32'd185;
#400 gamma=32'd1;row=32'd313;
#400 gamma=32'd5;row=32'd370;
#400 gamma=32'd1;row=32'd491;
#400 gamma=32'd4;row=32'd416;
#400 gamma=32'd2;row=32'd543;
#400 gamma=32'd2;row=32'd119;
#400 gamma=32'd2;row=32'd555;
#400 gamma=32'd1;row=32'd72;
#400 gamma=32'd2;row=32'd260;
#400 gamma=32'd3;row=32'd74;
#400 gamma=32'd1;row=32'd19;
#400 gamma=32'd3;row=32'd180;
#400 gamma=32'd3;row=32'd110;
#400 gamma=32'd4;row=32'd318;
#400 gamma=32'd1;row=32'd359;
#400 gamma=32'd5;row=32'd279;
#400 gamma=32'd4;row=32'd517;
#400 gamma=32'd5;row=32'd234;
#400 gamma=32'd5;row=32'd147;
#400 gamma=32'd4;row=32'd336;
#400 gamma=32'd4;row=32'd337;
#400 gamma=32'd1;row=32'd393;
#400 gamma=32'd1;row=32'd368;
#400 gamma=32'd1;row=32'd218;
#400 gamma=32'd4;row=32'd388;
#400 gamma=32'd1;row=32'd1;
#400 gamma=32'd3;row=32'd394;
#400 gamma=32'd2;row=32'd324;
#400 gamma=32'd3;row=32'd149;
#400 gamma=32'd5;row=32'd162;
#400 gamma=32'd4;row=32'd6;
#400 gamma=32'd4;row=32'd19;
#400 gamma=32'd4;row=32'd137;
#400 gamma=32'd4;row=32'd255;
#400 gamma=32'd5;row=32'd380;
#400 gamma=32'd5;row=32'd372;
#400 gamma=32'd1;row=32'd551;
#400 gamma=32'd1;row=32'd203;
#400 gamma=32'd4;row=32'd6;
#400 gamma=32'd3;row=32'd414;
#400 gamma=32'd1;row=32'd505;
#400 gamma=32'd1;row=32'd422;
#400 gamma=32'd3;row=32'd310;
#400 gamma=32'd5;row=32'd431;
#400 gamma=32'd3;row=32'd202;
#400 gamma=32'd2;row=32'd468;
#400 gamma=32'd4;row=32'd277;
#400 gamma=32'd4;row=32'd114;
#400 gamma=32'd1;row=32'd292;
#400 gamma=32'd5;row=32'd13;
#400 gamma=32'd4;row=32'd473;
#400 gamma=32'd3;row=32'd154;
#400 gamma=32'd2;row=32'd355;
#400 gamma=32'd5;row=32'd59;
#400 gamma=32'd5;row=32'd363;
#400 gamma=32'd5;row=32'd537;
#400 gamma=32'd3;row=32'd409;
#400 gamma=32'd5;row=32'd318;
#400 gamma=32'd5;row=32'd131;
#400 gamma=32'd2;row=32'd7;
#400 gamma=32'd1;row=32'd434;
#400 gamma=32'd1;row=32'd274;
#400 gamma=32'd5;row=32'd223;
#400 gamma=32'd4;row=32'd273;
#400 gamma=32'd2;row=32'd122;
#400 gamma=32'd2;row=32'd71;
#400 gamma=32'd2;row=32'd535;
#400 gamma=32'd4;row=32'd514;
#400 gamma=32'd5;row=32'd360;
#400 gamma=32'd3;row=32'd89;
#400 gamma=32'd5;row=32'd174;
#400 gamma=32'd5;row=32'd257;
#400 gamma=32'd3;row=32'd418;
#400 gamma=32'd3;row=32'd278;
#400 gamma=32'd1;row=32'd7;
#400 gamma=32'd4;row=32'd44;
#400 gamma=32'd1;row=32'd523;
#400 gamma=32'd3;row=32'd369;
#400 gamma=32'd4;row=32'd279;
#400 gamma=32'd5;row=32'd203;
#400 gamma=32'd2;row=32'd367;
#400 gamma=32'd2;row=32'd246;
#400 gamma=32'd1;row=32'd212;
#400 gamma=32'd4;row=32'd220;
#400 gamma=32'd1;row=32'd419;
#400 gamma=32'd4;row=32'd536;
#400 gamma=32'd2;row=32'd263;
#400 gamma=32'd5;row=32'd14;
#400 gamma=32'd1;row=32'd280;
#400 gamma=32'd5;row=32'd521;
#400 gamma=32'd3;row=32'd541;
#400 gamma=32'd1;row=32'd203;
#400 gamma=32'd4;row=32'd401;
#400 gamma=32'd2;row=32'd300;
#400 gamma=32'd3;row=32'd86;
#400 gamma=32'd2;row=32'd512;
#400 gamma=32'd1;row=32'd63;
#400 gamma=32'd3;row=32'd461;
#400 gamma=32'd4;row=32'd348;
#400 gamma=32'd3;row=32'd7;
#400 gamma=32'd5;row=32'd113;
#400 gamma=32'd3;row=32'd37;
#400 gamma=32'd4;row=32'd494;
#400 gamma=32'd2;row=32'd77;
#400 gamma=32'd1;row=32'd189;
#400 gamma=32'd2;row=32'd15;
#400 gamma=32'd1;row=32'd88;
#400 gamma=32'd3;row=32'd380;
#400 gamma=32'd5;row=32'd461;
#400 gamma=32'd3;row=32'd17;
#400 gamma=32'd4;row=32'd464;
#400 gamma=32'd5;row=32'd50;
#400 gamma=32'd2;row=32'd353;
#400 gamma=32'd3;row=32'd194;
#400 gamma=32'd2;row=32'd173;
#400 gamma=32'd3;row=32'd90;
#400 gamma=32'd4;row=32'd321;
#400 gamma=32'd1;row=32'd534;
#400 gamma=32'd5;row=32'd509;
#400 gamma=32'd1;row=32'd371;
#400 gamma=32'd4;row=32'd24;
#400 gamma=32'd3;row=32'd263;
#400 gamma=32'd4;row=32'd59;
#400 gamma=32'd1;row=32'd491;
#400 gamma=32'd1;row=32'd137;
#400 gamma=32'd1;row=32'd71;
#400 gamma=32'd2;row=32'd58;
#400 gamma=32'd4;row=32'd211;
#400 gamma=32'd4;row=32'd354;
#400 gamma=32'd5;row=32'd245;
#400 gamma=32'd2;row=32'd113;
#400 gamma=32'd1;row=32'd445;
#400 gamma=32'd2;row=32'd399;
#400 gamma=32'd2;row=32'd190;
#400 gamma=32'd3;row=32'd312;
#400 gamma=32'd3;row=32'd426;
#400 gamma=32'd5;row=32'd149;
#400 gamma=32'd1;row=32'd330;
#400 gamma=32'd3;row=32'd321;
#400 gamma=32'd1;row=32'd453;
#400 gamma=32'd1;row=32'd53;
#400 gamma=32'd2;row=32'd426;
#400 gamma=32'd4;row=32'd411;
#400 gamma=32'd2;row=32'd367;
#400 gamma=32'd4;row=32'd416;
#400 gamma=32'd4;row=32'd297;
#400 gamma=32'd2;row=32'd280;
#400 gamma=32'd3;row=32'd247;
#400 gamma=32'd5;row=32'd111;
#400 gamma=32'd2;row=32'd175;
#400 gamma=32'd2;row=32'd338;
#400 gamma=32'd1;row=32'd136;
#400 gamma=32'd1;row=32'd376;
#400 gamma=32'd1;row=32'd342;
#400 gamma=32'd5;row=32'd221;
#400 gamma=32'd2;row=32'd256;
#400 gamma=32'd2;row=32'd332;
#400 gamma=32'd4;row=32'd179;
#400 gamma=32'd2;row=32'd361;
#400 gamma=32'd4;row=32'd171;
#400 gamma=32'd3;row=32'd48;
#400 gamma=32'd2;row=32'd211;
#400 gamma=32'd5;row=32'd402;
#400 gamma=32'd3;row=32'd112;
#400 gamma=32'd1;row=32'd131;
#400 gamma=32'd1;row=32'd488;
#400 gamma=32'd4;row=32'd29;
#400 gamma=32'd4;row=32'd92;
#400 gamma=32'd1;row=32'd372;
#400 gamma=32'd5;row=32'd50;
#400 gamma=32'd5;row=32'd218;
#400 gamma=32'd1;row=32'd120;
#400 gamma=32'd1;row=32'd553;
#400 gamma=32'd5;row=32'd144;
#400 gamma=32'd2;row=32'd299;
#400 gamma=32'd1;row=32'd106;
#400 gamma=32'd4;row=32'd536;
#400 gamma=32'd1;row=32'd543;
#400 gamma=32'd3;row=32'd19;
#400 gamma=32'd1;row=32'd446;
#400 gamma=32'd3;row=32'd259;
#400 gamma=32'd4;row=32'd169;
#400 gamma=32'd3;row=32'd332;
#400 gamma=32'd5;row=32'd506;
#400 gamma=32'd5;row=32'd105;
#400 gamma=32'd4;row=32'd350;
#400 gamma=32'd5;row=32'd224;
#400 gamma=32'd5;row=32'd366;
#400 gamma=32'd1;row=32'd441;
#400 gamma=32'd2;row=32'd62;
#400 gamma=32'd1;row=32'd215;
#400 gamma=32'd1;row=32'd492;
#400 gamma=32'd2;row=32'd56;
#400 gamma=32'd3;row=32'd85;
#400 gamma=32'd2;row=32'd399;
#400 gamma=32'd4;row=32'd126;
#400 gamma=32'd4;row=32'd305;
#400 gamma=32'd2;row=32'd100;
#400 gamma=32'd1;row=32'd460;
#400 gamma=32'd2;row=32'd13;
#400 gamma=32'd5;row=32'd270;
#400 gamma=32'd2;row=32'd188;
#400 gamma=32'd2;row=32'd530;
#400 gamma=32'd5;row=32'd479;
#400 gamma=32'd1;row=32'd369;
#400 gamma=32'd2;row=32'd400;
#400 gamma=32'd5;row=32'd417;
#400 gamma=32'd2;row=32'd495;
#400 gamma=32'd2;row=32'd6;
#400 gamma=32'd4;row=32'd480;
#400 gamma=32'd3;row=32'd507;
#400 gamma=32'd5;row=32'd435;
#400 gamma=32'd4;row=32'd34;
#400 gamma=32'd5;row=32'd320;
#400 gamma=32'd1;row=32'd44;
#400 gamma=32'd4;row=32'd205;
#400 gamma=32'd3;row=32'd285;
#400 gamma=32'd5;row=32'd6;
#400 gamma=32'd4;row=32'd109;
#400 gamma=32'd1;row=32'd194;
#400 gamma=32'd1;row=32'd106;
#400 gamma=32'd1;row=32'd5;
#400 gamma=32'd4;row=32'd367;
#400 gamma=32'd2;row=32'd67;
#400 gamma=32'd4;row=32'd559;
#400 gamma=32'd4;row=32'd284;
#400 gamma=32'd4;row=32'd238;
#400 gamma=32'd5;row=32'd270;
#400 gamma=32'd4;row=32'd320;
#400 gamma=32'd1;row=32'd494;
#400 gamma=32'd2;row=32'd58;
#400 gamma=32'd5;row=32'd513;
#400 gamma=32'd2;row=32'd282;
#400 gamma=32'd5;row=32'd230;
#400 gamma=32'd4;row=32'd60;
#400 gamma=32'd4;row=32'd2;
#400 gamma=32'd5;row=32'd221;
#400 gamma=32'd3;row=32'd538;
#400 gamma=32'd5;row=32'd339;
#400 gamma=32'd2;row=32'd195;
#400 gamma=32'd5;row=32'd530;
#400 gamma=32'd1;row=32'd463;
#400 gamma=32'd2;row=32'd516;
#400 gamma=32'd2;row=32'd125;
#400 gamma=32'd1;row=32'd90;
#400 gamma=32'd1;row=32'd448;
#400 gamma=32'd4;row=32'd515;
#400 gamma=32'd1;row=32'd466;
#400 gamma=32'd1;row=32'd47;
#400 gamma=32'd1;row=32'd249;
#400 gamma=32'd5;row=32'd288;
#400 gamma=32'd4;row=32'd349;
#400 gamma=32'd5;row=32'd47;
#400 gamma=32'd4;row=32'd457;
#400 gamma=32'd3;row=32'd90;
#400 gamma=32'd2;row=32'd495;
#400 gamma=32'd3;row=32'd294;
#400 gamma=32'd4;row=32'd154;
#400 gamma=32'd3;row=32'd72;
#400 gamma=32'd4;row=32'd349;
#400 gamma=32'd1;row=32'd310;
#400 gamma=32'd2;row=32'd147;
#400 gamma=32'd1;row=32'd467;
#400 gamma=32'd3;row=32'd430;
#400 gamma=32'd4;row=32'd148;
#400 gamma=32'd2;row=32'd490;
#400 gamma=32'd2;row=32'd428;
#400 gamma=32'd5;row=32'd269;
#400 gamma=32'd3;row=32'd29;
#400 gamma=32'd4;row=32'd554;
#400 gamma=32'd2;row=32'd500;
#400 gamma=32'd4;row=32'd458;
#400 gamma=32'd3;row=32'd282;
#400 gamma=32'd1;row=32'd459;
#400 gamma=32'd1;row=32'd492;
#400 gamma=32'd2;row=32'd56;
#400 gamma=32'd4;row=32'd202;
#400 gamma=32'd4;row=32'd177;
#400 gamma=32'd5;row=32'd528;
#400 gamma=32'd2;row=32'd340;
#400 gamma=32'd2;row=32'd281;
#400 gamma=32'd3;row=32'd372;
#400 gamma=32'd2;row=32'd59;
#400 gamma=32'd1;row=32'd100;
#400 gamma=32'd2;row=32'd548;
#400 gamma=32'd3;row=32'd56;
#400 gamma=32'd5;row=32'd271;
#400 gamma=32'd2;row=32'd160;
#400 gamma=32'd5;row=32'd508;
#400 gamma=32'd4;row=32'd329;
#400 gamma=32'd1;row=32'd162;
#400 gamma=32'd2;row=32'd406;
#400 gamma=32'd5;row=32'd252;
#400 gamma=32'd2;row=32'd296;
#400 gamma=32'd3;row=32'd343;
#400 gamma=32'd3;row=32'd215;
#400 gamma=32'd1;row=32'd7;
#400 gamma=32'd3;row=32'd227;
#400 gamma=32'd2;row=32'd411;
#400 gamma=32'd3;row=32'd220;
#400 gamma=32'd5;row=32'd147;
#400 gamma=32'd4;row=32'd559;
#400 gamma=32'd5;row=32'd489;
#400 gamma=32'd5;row=32'd121;
#400 gamma=32'd1;row=32'd553;
#400 gamma=32'd2;row=32'd482;
#400 gamma=32'd3;row=32'd379;
#400 gamma=32'd2;row=32'd139;
#400 gamma=32'd5;row=32'd326;
#400 gamma=32'd4;row=32'd262;
#400 gamma=32'd2;row=32'd240;
#400 gamma=32'd4;row=32'd324;
#400 gamma=32'd5;row=32'd235;
#400 gamma=32'd2;row=32'd126;
#400 gamma=32'd5;row=32'd410;
#400 gamma=32'd1;row=32'd7;
#400 gamma=32'd3;row=32'd0;
#400 gamma=32'd2;row=32'd402;
#400 gamma=32'd1;row=32'd228;
#400 gamma=32'd5;row=32'd166;
#400 gamma=32'd3;row=32'd525;
#400 gamma=32'd2;row=32'd346;
#400 gamma=32'd1;row=32'd478;
#400 gamma=32'd1;row=32'd460;
#400 gamma=32'd2;row=32'd290;
#400 gamma=32'd1;row=32'd122;
#400 gamma=32'd3;row=32'd331;
#400 gamma=32'd4;row=32'd521;
#400 gamma=32'd2;row=32'd199;
#400 gamma=32'd2;row=32'd305;
#400 gamma=32'd5;row=32'd105;
#400 gamma=32'd4;row=32'd251;
#400 gamma=32'd2;row=32'd112;
#400 gamma=32'd3;row=32'd297;
#400 gamma=32'd5;row=32'd230;
#400 gamma=32'd4;row=32'd267;
#400 gamma=32'd3;row=32'd309;
#400 gamma=32'd3;row=32'd368;
#400 gamma=32'd1;row=32'd13;
#400 gamma=32'd2;row=32'd555;
#400 gamma=32'd3;row=32'd552;
#400 gamma=32'd2;row=32'd498;
#400 gamma=32'd1;row=32'd105;
#400 gamma=32'd5;row=32'd423;
#400 gamma=32'd2;row=32'd364;
#400 gamma=32'd5;row=32'd163;
#400 gamma=32'd5;row=32'd237;
#400 gamma=32'd4;row=32'd23;
#400 gamma=32'd5;row=32'd154;
#400 gamma=32'd5;row=32'd356;
#400 gamma=32'd4;row=32'd382;
#400 gamma=32'd3;row=32'd263;
#400 gamma=32'd5;row=32'd32;
#400 gamma=32'd3;row=32'd379;
#400 gamma=32'd3;row=32'd113;
#400 gamma=32'd5;row=32'd387;
#400 gamma=32'd3;row=32'd4;
#400 gamma=32'd4;row=32'd448;
#400 gamma=32'd3;row=32'd413;
#400 gamma=32'd3;row=32'd512;
#400 gamma=32'd2;row=32'd546;
#400 gamma=32'd1;row=32'd268;
#400 gamma=32'd4;row=32'd510;
#400 gamma=32'd4;row=32'd57;
#400 gamma=32'd3;row=32'd395;
#400 gamma=32'd1;row=32'd89;
#400 gamma=32'd4;row=32'd469;
#400 gamma=32'd4;row=32'd496;
#400 gamma=32'd1;row=32'd273;
#400 gamma=32'd5;row=32'd479;
#400 gamma=32'd4;row=32'd446;
#400 gamma=32'd1;row=32'd33;
#400 gamma=32'd2;row=32'd327;
#400 gamma=32'd1;row=32'd48;
#400 gamma=32'd4;row=32'd517;
#400 gamma=32'd5;row=32'd522;
#400 gamma=32'd2;row=32'd92;
#400 gamma=32'd4;row=32'd535;
#400 gamma=32'd5;row=32'd465;
#400 gamma=32'd3;row=32'd558;
#400 gamma=32'd3;row=32'd237;
#400 gamma=32'd2;row=32'd438;
#400 gamma=32'd4;row=32'd122;
#400 gamma=32'd5;row=32'd199;
#400 gamma=32'd1;row=32'd255;
#400 gamma=32'd1;row=32'd59;
#400 gamma=32'd3;row=32'd550;
#400 gamma=32'd4;row=32'd538;
#400 gamma=32'd5;row=32'd99;
#400 gamma=32'd4;row=32'd38;
#400 gamma=32'd2;row=32'd75;
#400 gamma=32'd4;row=32'd330;
#400 gamma=32'd5;row=32'd209;
#400 gamma=32'd5;row=32'd245;
#400 gamma=32'd1;row=32'd157;
#400 gamma=32'd1;row=32'd342;
#400 gamma=32'd1;row=32'd266;
#400 gamma=32'd1;row=32'd318;
#400 gamma=32'd2;row=32'd275;
#400 gamma=32'd2;row=32'd310;
#400 gamma=32'd3;row=32'd198;
#400 gamma=32'd4;row=32'd150;
#400 gamma=32'd2;row=32'd430;
#400 gamma=32'd1;row=32'd311;
#400 gamma=32'd2;row=32'd98;
#400 gamma=32'd2;row=32'd475;
#400 gamma=32'd5;row=32'd103;
#400 gamma=32'd1;row=32'd445;
#400 gamma=32'd3;row=32'd18;
#400 gamma=32'd4;row=32'd469;
#400 gamma=32'd3;row=32'd67;
#400 gamma=32'd5;row=32'd211;
#400 gamma=32'd4;row=32'd112;
#400 gamma=32'd3;row=32'd110;
#400 gamma=32'd2;row=32'd48;
#400 gamma=32'd5;row=32'd51;
#400 gamma=32'd5;row=32'd115;
#400 gamma=32'd1;row=32'd227;
#400 gamma=32'd5;row=32'd280;
#400 gamma=32'd5;row=32'd100;
#400 gamma=32'd2;row=32'd113;
#400 gamma=32'd3;row=32'd412;
#400 gamma=32'd3;row=32'd542;
#400 gamma=32'd3;row=32'd527;
#400 gamma=32'd1;row=32'd48;
#400 gamma=32'd2;row=32'd262;
#400 gamma=32'd4;row=32'd549;
#400 gamma=32'd1;row=32'd390;
#400 gamma=32'd5;row=32'd327;
#400 gamma=32'd1;row=32'd506;
#400 gamma=32'd1;row=32'd410;
#400 gamma=32'd5;row=32'd513;
#400 gamma=32'd2;row=32'd121;
#400 gamma=32'd3;row=32'd325;
#400 gamma=32'd2;row=32'd441;
#400 gamma=32'd4;row=32'd25;
#400 gamma=32'd4;row=32'd337;
#400 gamma=32'd2;row=32'd110;
#400 gamma=32'd4;row=32'd409;
#400 gamma=32'd2;row=32'd74;
#400 gamma=32'd2;row=32'd127;
#400 gamma=32'd1;row=32'd474;
#400 gamma=32'd5;row=32'd200;
#400 gamma=32'd3;row=32'd107;
#400 gamma=32'd4;row=32'd539;
#400 gamma=32'd4;row=32'd158;
#400 gamma=32'd4;row=32'd149;
#400 gamma=32'd1;row=32'd239;
#400 gamma=32'd3;row=32'd305;
#400 gamma=32'd4;row=32'd282;
#400 gamma=32'd1;row=32'd391;
#400 gamma=32'd3;row=32'd276;
#400 gamma=32'd4;row=32'd193;
#400 gamma=32'd2;row=32'd552;
#400 gamma=32'd2;row=32'd26;
#400 gamma=32'd4;row=32'd189;
#400 gamma=32'd1;row=32'd437;
#400 gamma=32'd2;row=32'd217;
#400 gamma=32'd3;row=32'd503;
#400 gamma=32'd3;row=32'd107;
#400 gamma=32'd3;row=32'd469;
#400 gamma=32'd1;row=32'd445;
#400 gamma=32'd2;row=32'd231;
#400 gamma=32'd5;row=32'd108;
#400 gamma=32'd5;row=32'd150;
#400 gamma=32'd1;row=32'd107;
#400 gamma=32'd1;row=32'd244;
#400 gamma=32'd2;row=32'd356;
#400 gamma=32'd1;row=32'd396;
#400 gamma=32'd1;row=32'd375;
#400 gamma=32'd5;row=32'd363;
#400 gamma=32'd3;row=32'd284;
#400 gamma=32'd2;row=32'd351;
#400 gamma=32'd2;row=32'd510;
#400 gamma=32'd1;row=32'd400;
#400 gamma=32'd5;row=32'd51;
#400 gamma=32'd1;row=32'd422;
#400 gamma=32'd1;row=32'd48;
#400 gamma=32'd2;row=32'd215;
#400 gamma=32'd1;row=32'd324;
#400 gamma=32'd5;row=32'd50;
#400 gamma=32'd1;row=32'd438;
#400 gamma=32'd2;row=32'd378;
#400 gamma=32'd4;row=32'd86;
#400 gamma=32'd2;row=32'd423;
#400 gamma=32'd3;row=32'd16;
#400 gamma=32'd5;row=32'd169;
#400 gamma=32'd5;row=32'd195;
#400 gamma=32'd4;row=32'd301;
#400 gamma=32'd2;row=32'd460;
#400 gamma=32'd2;row=32'd293;
#400 gamma=32'd1;row=32'd260;
#400 gamma=32'd4;row=32'd550;
#400 gamma=32'd5;row=32'd511;
#400 gamma=32'd5;row=32'd504;
#400 gamma=32'd5;row=32'd407;
#400 gamma=32'd4;row=32'd483;
#400 gamma=32'd5;row=32'd238;
#400 gamma=32'd5;row=32'd21;
#400 gamma=32'd3;row=32'd462;
#400 gamma=32'd5;row=32'd343;
#400 gamma=32'd2;row=32'd249;
#400 gamma=32'd5;row=32'd57;
#400 gamma=32'd4;row=32'd270;
#400 gamma=32'd5;row=32'd268;
#400 gamma=32'd2;row=32'd559;
#400 gamma=32'd5;row=32'd424;
#400 gamma=32'd1;row=32'd359;
#400 gamma=32'd5;row=32'd390;
#400 gamma=32'd5;row=32'd32;
#400 gamma=32'd1;row=32'd56;
#400 gamma=32'd5;row=32'd526;
#400 gamma=32'd2;row=32'd547;
#400 gamma=32'd2;row=32'd420;
#400 gamma=32'd1;row=32'd149;
#400 gamma=32'd4;row=32'd452;
#400 gamma=32'd1;row=32'd434;
#400 gamma=32'd3;row=32'd284;
#400 gamma=32'd1;row=32'd477;
#400 gamma=32'd1;row=32'd57;
#400 gamma=32'd5;row=32'd352;
#400 gamma=32'd5;row=32'd190;
#400 gamma=32'd4;row=32'd555;
#400 gamma=32'd5;row=32'd250;
#400 gamma=32'd3;row=32'd28;
#400 gamma=32'd3;row=32'd105;
#400 gamma=32'd3;row=32'd447;
#400 gamma=32'd2;row=32'd184;
#400 gamma=32'd1;row=32'd419;
#400 gamma=32'd2;row=32'd427;
#400 gamma=32'd3;row=32'd498;
#400 gamma=32'd3;row=32'd363;
#400 gamma=32'd5;row=32'd151;
#400 gamma=32'd5;row=32'd219;
#400 gamma=32'd1;row=32'd434;
#400 gamma=32'd5;row=32'd398;
#400 gamma=32'd4;row=32'd522;
#400 gamma=32'd2;row=32'd333;
#400 gamma=32'd3;row=32'd110;
#400 gamma=32'd5;row=32'd188;
#400 gamma=32'd5;row=32'd285;
#400 gamma=32'd5;row=32'd325;
#400 gamma=32'd2;row=32'd202;
#400 gamma=32'd3;row=32'd186;
#400 gamma=32'd2;row=32'd431;
#400 gamma=32'd4;row=32'd108;
#400 gamma=32'd1;row=32'd374;
#400 gamma=32'd4;row=32'd132;
#400 gamma=32'd4;row=32'd84;
#400 gamma=32'd3;row=32'd195;
#400 gamma=32'd3;row=32'd80;
#400 gamma=32'd1;row=32'd160;
#400 gamma=32'd5;row=32'd156;
#400 gamma=32'd3;row=32'd508;
#400 gamma=32'd5;row=32'd277;
#400 gamma=32'd4;row=32'd229;
#400 gamma=32'd4;row=32'd511;
#400 gamma=32'd1;row=32'd128;
#400 gamma=32'd2;row=32'd277;
#400 gamma=32'd2;row=32'd144;
#400 gamma=32'd4;row=32'd486;
#400 gamma=32'd2;row=32'd265;
#400 gamma=32'd1;row=32'd116;
#400 gamma=32'd5;row=32'd102;
#400 gamma=32'd1;row=32'd16;
#400 gamma=32'd4;row=32'd158;
#400 gamma=32'd5;row=32'd71;
#400 gamma=32'd5;row=32'd479;
#400 gamma=32'd1;row=32'd144;
#400 gamma=32'd4;row=32'd88;
#400 gamma=32'd5;row=32'd170;
#400 gamma=32'd3;row=32'd42;
#400 gamma=32'd2;row=32'd444;
#400 gamma=32'd1;row=32'd472;
#400 gamma=32'd3;row=32'd291;
#400 gamma=32'd3;row=32'd37;
#400 gamma=32'd2;row=32'd199;
#400 gamma=32'd4;row=32'd183;
#400 gamma=32'd2;row=32'd62;
#400 gamma=32'd1;row=32'd283;
#400 gamma=32'd3;row=32'd444;
#400 gamma=32'd2;row=32'd227;
#400 gamma=32'd3;row=32'd253;
#400 gamma=32'd4;row=32'd198;
#400 gamma=32'd3;row=32'd425;
#400 gamma=32'd4;row=32'd171;
#400 gamma=32'd1;row=32'd412;
#400 gamma=32'd1;row=32'd385;
#400 gamma=32'd4;row=32'd351;
#400 gamma=32'd5;row=32'd212;
#400 gamma=32'd5;row=32'd262;
#400 gamma=32'd2;row=32'd268;
#400 gamma=32'd4;row=32'd147;
#400 gamma=32'd3;row=32'd1;
#400 gamma=32'd5;row=32'd356;
#400 gamma=32'd1;row=32'd66;
#400 gamma=32'd1;row=32'd75;
#400 gamma=32'd4;row=32'd388;
#400 gamma=32'd2;row=32'd285;
#400 gamma=32'd5;row=32'd62;
#400 gamma=32'd4;row=32'd172;
#400 gamma=32'd2;row=32'd322;
#400 gamma=32'd5;row=32'd293;
#400 gamma=32'd4;row=32'd376;
#400 gamma=32'd2;row=32'd427;
#400 gamma=32'd1;row=32'd426;
#400 gamma=32'd3;row=32'd85;
#400 gamma=32'd2;row=32'd318;
#400 gamma=32'd1;row=32'd290;
#400 gamma=32'd1;row=32'd266;
#400 gamma=32'd5;row=32'd13;
#400 gamma=32'd1;row=32'd372;
#400 gamma=32'd3;row=32'd198;
#400 gamma=32'd1;row=32'd517;
#400 gamma=32'd2;row=32'd462;
#400 gamma=32'd5;row=32'd93;
#400 gamma=32'd3;row=32'd114;
#400 gamma=32'd5;row=32'd35;
#400 gamma=32'd1;row=32'd173;
#400 gamma=32'd5;row=32'd229;
#400 gamma=32'd4;row=32'd115;
#400 gamma=32'd2;row=32'd391;
#400 gamma=32'd4;row=32'd239;
#400 gamma=32'd4;row=32'd384;
#400 gamma=32'd3;row=32'd275;
#400 gamma=32'd1;row=32'd285;
#400 gamma=32'd1;row=32'd89;
#400 gamma=32'd3;row=32'd78;
#400 gamma=32'd2;row=32'd293;
#400 gamma=32'd4;row=32'd88;
#400 gamma=32'd3;row=32'd320;
#400 gamma=32'd2;row=32'd63;
#400 gamma=32'd2;row=32'd281;
#400 gamma=32'd3;row=32'd403;
#400 gamma=32'd5;row=32'd377;
#400 gamma=32'd3;row=32'd447;
#400 gamma=32'd2;row=32'd61;
#400 gamma=32'd2;row=32'd344;
#400 gamma=32'd4;row=32'd530;
#400 gamma=32'd5;row=32'd355;
#400 gamma=32'd3;row=32'd91;
#400 gamma=32'd5;row=32'd533;
#400 gamma=32'd4;row=32'd422;
#400 gamma=32'd2;row=32'd431;
#400 gamma=32'd4;row=32'd534;
#400 gamma=32'd3;row=32'd148;
#400 gamma=32'd5;row=32'd389;
#400 gamma=32'd4;row=32'd540;
#400 gamma=32'd3;row=32'd332;
#400 gamma=32'd2;row=32'd37;
#400 gamma=32'd1;row=32'd519;
#400 gamma=32'd1;row=32'd240;
#400 gamma=32'd1;row=32'd165;
#400 gamma=32'd2;row=32'd184;
#400 gamma=32'd1;row=32'd99;
#400 gamma=32'd2;row=32'd71;
#400 gamma=32'd5;row=32'd2;
#400 gamma=32'd3;row=32'd162;
#400 gamma=32'd1;row=32'd108;
#400 gamma=32'd4;row=32'd454;
#400 gamma=32'd2;row=32'd86;
#400 gamma=32'd3;row=32'd62;
#400 gamma=32'd3;row=32'd142;
#400 gamma=32'd5;row=32'd429;
#400 gamma=32'd5;row=32'd511;
#400 gamma=32'd3;row=32'd454;
#400 gamma=32'd4;row=32'd38;
#400 gamma=32'd5;row=32'd101;
#400 gamma=32'd1;row=32'd518;
#400 gamma=32'd1;row=32'd11;
#400 gamma=32'd5;row=32'd308;
#400 gamma=32'd5;row=32'd524;
#400 gamma=32'd4;row=32'd8;
#400 gamma=32'd1;row=32'd141;
#400 gamma=32'd1;row=32'd404;
#400 gamma=32'd1;row=32'd393;
#400 gamma=32'd2;row=32'd345;
#400 gamma=32'd5;row=32'd290;
#400 gamma=32'd3;row=32'd184;
#400 gamma=32'd4;row=32'd85;
#400 gamma=32'd2;row=32'd486;
#400 gamma=32'd5;row=32'd513;
#400 gamma=32'd3;row=32'd504;
#400 gamma=32'd1;row=32'd415;
#400 gamma=32'd4;row=32'd281;
#400 gamma=32'd4;row=32'd118;
#400 gamma=32'd5;row=32'd136;
#400 gamma=32'd1;row=32'd446;
#400 gamma=32'd4;row=32'd35;
#400 gamma=32'd5;row=32'd6;
#400 gamma=32'd2;row=32'd170;
#400 gamma=32'd5;row=32'd301;
#400 gamma=32'd1;row=32'd448;
#400 gamma=32'd4;row=32'd54;
#400 gamma=32'd4;row=32'd410;
#400 gamma=32'd4;row=32'd55;
#400 gamma=32'd1;row=32'd507;
#400 gamma=32'd2;row=32'd503;
#400 gamma=32'd3;row=32'd518;
#400 gamma=32'd3;row=32'd46;
#400 gamma=32'd4;row=32'd349;
#400 gamma=32'd5;row=32'd451;
#400 gamma=32'd3;row=32'd227;
#400 gamma=32'd1;row=32'd107;
#400 gamma=32'd4;row=32'd228;
#400 gamma=32'd1;row=32'd448;
#400 gamma=32'd2;row=32'd42;
#400 gamma=32'd3;row=32'd101;
#400 gamma=32'd3;row=32'd390;
#400 gamma=32'd1;row=32'd174;
#400 gamma=32'd5;row=32'd0;
#400 gamma=32'd5;row=32'd436;
#400 gamma=32'd5;row=32'd141;
#400 gamma=32'd3;row=32'd433;
#400 gamma=32'd4;row=32'd96;
#400 gamma=32'd5;row=32'd186;
#400 gamma=32'd3;row=32'd136;
#400 gamma=32'd2;row=32'd141;
#400 gamma=32'd5;row=32'd238;
#400 gamma=32'd4;row=32'd265;
#400 gamma=32'd5;row=32'd496;
#400 gamma=32'd1;row=32'd328;
#400 gamma=32'd1;row=32'd124;
#400 gamma=32'd4;row=32'd374;
#400 gamma=32'd5;row=32'd157;
#400 gamma=32'd5;row=32'd199;
#400 gamma=32'd1;row=32'd404;
#400 gamma=32'd3;row=32'd472;
#400 gamma=32'd5;row=32'd89;
#400 gamma=32'd5;row=32'd35;
#400 gamma=32'd5;row=32'd178;
#400 gamma=32'd1;row=32'd536;
#400 gamma=32'd3;row=32'd452;
#400 gamma=32'd4;row=32'd400;
#400 gamma=32'd2;row=32'd271;
#400 gamma=32'd2;row=32'd114;
#400 gamma=32'd5;row=32'd189;
#400 gamma=32'd1;row=32'd151;
#400 gamma=32'd1;row=32'd241;
#400 gamma=32'd5;row=32'd63;
#400 gamma=32'd4;row=32'd131;
#400 gamma=32'd5;row=32'd246;
#400 gamma=32'd5;row=32'd265;
#400 gamma=32'd3;row=32'd142;
#400 gamma=32'd1;row=32'd170;
#400 gamma=32'd1;row=32'd356;
#400 gamma=32'd2;row=32'd541;
#400 gamma=32'd2;row=32'd206;
#400 gamma=32'd3;row=32'd162;
#400 gamma=32'd4;row=32'd508;
#400 gamma=32'd3;row=32'd20;
#400 gamma=32'd5;row=32'd406;
#400 gamma=32'd1;row=32'd552;
#400 gamma=32'd5;row=32'd500;
#400 gamma=32'd5;row=32'd136;
#400 gamma=32'd4;row=32'd339;
#400 gamma=32'd1;row=32'd40;
#400 gamma=32'd2;row=32'd279;
#400 gamma=32'd4;row=32'd262;
#400 gamma=32'd2;row=32'd289;
#400 gamma=32'd5;row=32'd318;
#400 gamma=32'd1;row=32'd552;
#400 gamma=32'd3;row=32'd71;
#400 gamma=32'd5;row=32'd38;
#400 gamma=32'd3;row=32'd415;
#400 gamma=32'd2;row=32'd410;
#400 gamma=32'd2;row=32'd170;
#400 gamma=32'd5;row=32'd543;
#400 gamma=32'd5;row=32'd313;
#400 gamma=32'd2;row=32'd338;
#400 gamma=32'd3;row=32'd174;
#400 gamma=32'd5;row=32'd320;
#400 gamma=32'd5;row=32'd163;
#400 gamma=32'd1;row=32'd252;
#400 gamma=32'd5;row=32'd344;
#400 gamma=32'd4;row=32'd407;
#400 gamma=32'd4;row=32'd102;
#400 gamma=32'd1;row=32'd414;
#400 gamma=32'd1;row=32'd34;
#400 gamma=32'd5;row=32'd374;
#400 gamma=32'd1;row=32'd522;
#400 gamma=32'd1;row=32'd415;
#400 gamma=32'd3;row=32'd364;
#400 gamma=32'd4;row=32'd206;
#400 gamma=32'd1;row=32'd241;
#400 gamma=32'd4;row=32'd267;
#400 gamma=32'd5;row=32'd378;
#400 gamma=32'd5;row=32'd301;
#400 gamma=32'd5;row=32'd158;
#400 gamma=32'd1;row=32'd224;
#400 gamma=32'd3;row=32'd316;
#400 gamma=32'd4;row=32'd451;
#400 gamma=32'd5;row=32'd319;
#400 gamma=32'd2;row=32'd383;
#400 gamma=32'd4;row=32'd494;
#400 gamma=32'd1;row=32'd488;
#400 gamma=32'd5;row=32'd368;
#400 gamma=32'd1;row=32'd421;
#400 gamma=32'd5;row=32'd234;
#400 gamma=32'd3;row=32'd422;
#400 gamma=32'd1;row=32'd298;
#400 gamma=32'd3;row=32'd138;
#400 gamma=32'd2;row=32'd556;
#400 gamma=32'd5;row=32'd135;
#400 gamma=32'd2;row=32'd25;
#400 gamma=32'd3;row=32'd209;
#400 gamma=32'd5;row=32'd474;
#400 gamma=32'd5;row=32'd477;
#400 gamma=32'd3;row=32'd522;
#400 gamma=32'd1;row=32'd42;
#400 gamma=32'd1;row=32'd70;
#400 gamma=32'd4;row=32'd417;
#400 gamma=32'd3;row=32'd239;
#400 gamma=32'd3;row=32'd95;
#400 gamma=32'd1;row=32'd44;
#400 gamma=32'd2;row=32'd133;
#400 gamma=32'd1;row=32'd48;
#400 gamma=32'd2;row=32'd433;
#400 gamma=32'd5;row=32'd27;
#400 gamma=32'd4;row=32'd106;
#400 gamma=32'd3;row=32'd135;
#400 gamma=32'd5;row=32'd356;
#400 gamma=32'd3;row=32'd435;
#400 gamma=32'd1;row=32'd211;
#400 gamma=32'd2;row=32'd385;
#400 gamma=32'd1;row=32'd525;
#400 gamma=32'd2;row=32'd257;
#400 gamma=32'd2;row=32'd72;
#400 gamma=32'd2;row=32'd129;
#400 gamma=32'd1;row=32'd103;
#400 gamma=32'd2;row=32'd407;
#400 gamma=32'd2;row=32'd68;
#400 gamma=32'd3;row=32'd443;
#400 gamma=32'd4;row=32'd279;
#400 gamma=32'd3;row=32'd195;
#400 gamma=32'd5;row=32'd169;
#400 gamma=32'd4;row=32'd185;
#400 gamma=32'd4;row=32'd201;
#400 gamma=32'd3;row=32'd73;
#400 gamma=32'd1;row=32'd323;
#400 gamma=32'd3;row=32'd351;
#400 gamma=32'd2;row=32'd111;
#400 gamma=32'd3;row=32'd312;
#400 gamma=32'd5;row=32'd510;
#400 gamma=32'd2;row=32'd475;
#400 gamma=32'd1;row=32'd163;
#400 gamma=32'd3;row=32'd279;
#400 gamma=32'd1;row=32'd111;
#400 gamma=32'd1;row=32'd133;
#400 gamma=32'd1;row=32'd289;
#400 gamma=32'd1;row=32'd142;
#400 gamma=32'd3;row=32'd471;
#400 gamma=32'd5;row=32'd60;
#400 gamma=32'd5;row=32'd430;
#400 gamma=32'd3;row=32'd51;
#400 gamma=32'd1;row=32'd516;
#400 gamma=32'd3;row=32'd59;
#400 gamma=32'd3;row=32'd261;
#400 gamma=32'd2;row=32'd38;
#400 gamma=32'd3;row=32'd158;
#400 gamma=32'd1;row=32'd162;
#400 gamma=32'd4;row=32'd490;
#400 gamma=32'd2;row=32'd121;
#400 gamma=32'd1;row=32'd315;
#400 gamma=32'd4;row=32'd412;
#400 gamma=32'd1;row=32'd392;
#400 gamma=32'd2;row=32'd304;
#400 gamma=32'd4;row=32'd310;
#400 gamma=32'd2;row=32'd220;
#400 gamma=32'd2;row=32'd390;
#400 gamma=32'd2;row=32'd310;
#400 gamma=32'd3;row=32'd274;
#400 gamma=32'd3;row=32'd279;
#400 gamma=32'd4;row=32'd454;
#400 gamma=32'd4;row=32'd154;
#400 gamma=32'd1;row=32'd137;
#400 gamma=32'd3;row=32'd238;
#400 gamma=32'd2;row=32'd288;
#400 gamma=32'd1;row=32'd329;
#400 gamma=32'd1;row=32'd89;
#400 gamma=32'd5;row=32'd488;
#400 gamma=32'd5;row=32'd212;
#400 gamma=32'd4;row=32'd314;
#400 gamma=32'd5;row=32'd527;
#400 gamma=32'd2;row=32'd256;
#400 gamma=32'd5;row=32'd26;
#400 gamma=32'd4;row=32'd348;
#400 gamma=32'd3;row=32'd167;
#400 gamma=32'd2;row=32'd400;
#400 gamma=32'd2;row=32'd247;
#400 gamma=32'd5;row=32'd383;
#400 gamma=32'd1;row=32'd511;
#400 gamma=32'd3;row=32'd136;
#400 gamma=32'd5;row=32'd526;
#400 gamma=32'd1;row=32'd524;
#400 gamma=32'd4;row=32'd541;
#400 gamma=32'd3;row=32'd26;
#400 gamma=32'd4;row=32'd327;
#400 gamma=32'd4;row=32'd378;
#400 gamma=32'd1;row=32'd202;
#400 gamma=32'd1;row=32'd425;
#400 gamma=32'd3;row=32'd235;
#400 gamma=32'd3;row=32'd293;
#400 gamma=32'd4;row=32'd205;
#400 gamma=32'd4;row=32'd347;
#400 gamma=32'd3;row=32'd356;
#400 gamma=32'd1;row=32'd125;
#400 gamma=32'd3;row=32'd340;
#400 gamma=32'd4;row=32'd56;
#400 gamma=32'd3;row=32'd91;
#400 gamma=32'd3;row=32'd470;
#400 gamma=32'd5;row=32'd501;
#400 gamma=32'd1;row=32'd304;
#400 gamma=32'd2;row=32'd548;
#400 gamma=32'd5;row=32'd61;
#400 gamma=32'd4;row=32'd267;
#400 gamma=32'd3;row=32'd444;
#400 gamma=32'd3;row=32'd306;
#400 gamma=32'd4;row=32'd218;
#400 gamma=32'd5;row=32'd114;
#400 gamma=32'd1;row=32'd170;
#400 gamma=32'd1;row=32'd30;
#400 gamma=32'd2;row=32'd500;
#400 gamma=32'd5;row=32'd396;
#400 gamma=32'd2;row=32'd66;
#400 gamma=32'd1;row=32'd482;
#400 gamma=32'd4;row=32'd158;
#400 gamma=32'd5;row=32'd558;
#400 gamma=32'd4;row=32'd495;
#400 gamma=32'd5;row=32'd290;
#400 gamma=32'd1;row=32'd283;
#400 gamma=32'd5;row=32'd553;
#400 gamma=32'd3;row=32'd204;
#400 gamma=32'd4;row=32'd159;
#400 gamma=32'd1;row=32'd392;
#400 gamma=32'd2;row=32'd458;
#400 gamma=32'd4;row=32'd513;
#400 gamma=32'd2;row=32'd213;
#400 gamma=32'd5;row=32'd481;
#400 gamma=32'd4;row=32'd243;
#400 gamma=32'd4;row=32'd25;
#400 gamma=32'd3;row=32'd129;
#400 gamma=32'd4;row=32'd557;
#400 gamma=32'd1;row=32'd284;
#400 gamma=32'd3;row=32'd324;
#400 gamma=32'd1;row=32'd255;
#400 gamma=32'd4;row=32'd218;
#400 gamma=32'd2;row=32'd236;
#400 gamma=32'd1;row=32'd95;
#400 gamma=32'd3;row=32'd104;
#400 gamma=32'd5;row=32'd287;
#400 gamma=32'd1;row=32'd489;
#400 gamma=32'd1;row=32'd372;
#400 gamma=32'd2;row=32'd81;
#400 gamma=32'd2;row=32'd22;
#400 gamma=32'd4;row=32'd362;
#400 gamma=32'd1;row=32'd268;
#400 gamma=32'd3;row=32'd11;
#400 gamma=32'd5;row=32'd268;
#400 gamma=32'd2;row=32'd360;
#400 gamma=32'd5;row=32'd371;
#400 gamma=32'd5;row=32'd381;
#400 gamma=32'd1;row=32'd559;
#400 gamma=32'd1;row=32'd153;
#400 gamma=32'd1;row=32'd54;
#400 gamma=32'd2;row=32'd196;
#400 gamma=32'd3;row=32'd526;
#400 gamma=32'd4;row=32'd518;
#400 gamma=32'd1;row=32'd41;
#400 gamma=32'd2;row=32'd154;
#400 gamma=32'd1;row=32'd7;
#400 gamma=32'd2;row=32'd285;
#400 gamma=32'd5;row=32'd218;
#400 gamma=32'd5;row=32'd70;
#400 gamma=32'd1;row=32'd324;
#400 gamma=32'd4;row=32'd80;
#400 gamma=32'd4;row=32'd104;
#400 gamma=32'd1;row=32'd44;
#400 gamma=32'd2;row=32'd77;
#400 gamma=32'd2;row=32'd396;
#400 gamma=32'd1;row=32'd272;
#400 gamma=32'd1;row=32'd350;
#400 gamma=32'd4;row=32'd208;
#400 gamma=32'd2;row=32'd299;
#400 gamma=32'd3;row=32'd29;
#400 gamma=32'd1;row=32'd435;
#400 gamma=32'd2;row=32'd380;
#400 gamma=32'd5;row=32'd551;
#400 gamma=32'd5;row=32'd439;
#400 gamma=32'd2;row=32'd191;
#400 gamma=32'd4;row=32'd274;
#400 gamma=32'd3;row=32'd426;
#400 gamma=32'd5;row=32'd42;
#400 gamma=32'd2;row=32'd160;
#400 gamma=32'd4;row=32'd1;
#400 gamma=32'd2;row=32'd9;
#400 gamma=32'd3;row=32'd432;
#400 gamma=32'd1;row=32'd295;
#400 gamma=32'd3;row=32'd87;
#400 gamma=32'd5;row=32'd60;
#400 gamma=32'd4;row=32'd87;
#400 gamma=32'd2;row=32'd301;
#400 gamma=32'd5;row=32'd215;
#400 gamma=32'd3;row=32'd137;
#400 gamma=32'd4;row=32'd48;
#400 gamma=32'd5;row=32'd211;
#400 gamma=32'd3;row=32'd114;
#400 gamma=32'd5;row=32'd504;
#400 gamma=32'd2;row=32'd248;
#400 gamma=32'd5;row=32'd127;
#400 gamma=32'd1;row=32'd85;
#400 gamma=32'd4;row=32'd224;
#400 gamma=32'd4;row=32'd392;
#400 gamma=32'd1;row=32'd491;
#400 gamma=32'd5;row=32'd428;
#400 gamma=32'd4;row=32'd19;
#400 gamma=32'd4;row=32'd375;
#400 gamma=32'd3;row=32'd269;
#400 gamma=32'd1;row=32'd57;
#400 gamma=32'd4;row=32'd189;
#400 gamma=32'd2;row=32'd359;
#400 gamma=32'd3;row=32'd21;
#400 gamma=32'd5;row=32'd209;
#400 gamma=32'd2;row=32'd433;
#400 gamma=32'd2;row=32'd522;
#400 gamma=32'd3;row=32'd498;
#400 gamma=32'd5;row=32'd280;
#400 gamma=32'd2;row=32'd533;
#400 gamma=32'd3;row=32'd483;
#400 gamma=32'd5;row=32'd293;
#400 gamma=32'd3;row=32'd202;
#400 gamma=32'd4;row=32'd290;
#400 gamma=32'd2;row=32'd176;
#400 gamma=32'd4;row=32'd170;
#400 gamma=32'd5;row=32'd115;
#400 gamma=32'd2;row=32'd13;
#400 gamma=32'd3;row=32'd26;
#400 gamma=32'd3;row=32'd478;
#400 gamma=32'd1;row=32'd475;
#400 gamma=32'd3;row=32'd442;
#400 gamma=32'd2;row=32'd401;
#400 gamma=32'd5;row=32'd318;
#400 gamma=32'd4;row=32'd46;
#400 gamma=32'd1;row=32'd167;
#400 gamma=32'd2;row=32'd432;
#400 gamma=32'd4;row=32'd330;
#400 gamma=32'd4;row=32'd306;
#400 gamma=32'd1;row=32'd466;
#400 gamma=32'd2;row=32'd254;
#400 gamma=32'd2;row=32'd511;
#400 gamma=32'd3;row=32'd56;
#400 gamma=32'd3;row=32'd243;
#400 gamma=32'd3;row=32'd99;
#400 gamma=32'd4;row=32'd233;
#400 gamma=32'd2;row=32'd205;
#400 gamma=32'd2;row=32'd42;
#400 gamma=32'd1;row=32'd301;
#400 gamma=32'd1;row=32'd208;
#400 gamma=32'd3;row=32'd153;
#400 gamma=32'd3;row=32'd334;
#400 gamma=32'd4;row=32'd219;
#400 gamma=32'd5;row=32'd419;
#400 gamma=32'd5;row=32'd330;
#400 gamma=32'd2;row=32'd87;
#400 gamma=32'd2;row=32'd416;
#400 gamma=32'd4;row=32'd512;
#400 gamma=32'd1;row=32'd47;
#400 gamma=32'd5;row=32'd305;
#400 gamma=32'd2;row=32'd11;
#400 gamma=32'd5;row=32'd399;
#400 gamma=32'd1;row=32'd528;
#400 gamma=32'd3;row=32'd198;
#400 gamma=32'd1;row=32'd303;
#400 gamma=32'd1;row=32'd62;
#400 gamma=32'd2;row=32'd92;
#400 gamma=32'd3;row=32'd146;
#400 gamma=32'd4;row=32'd552;
#400 gamma=32'd2;row=32'd89;
#400 gamma=32'd5;row=32'd49;
#400 gamma=32'd1;row=32'd332;
#400 gamma=32'd1;row=32'd178;
#400 gamma=32'd2;row=32'd356;
#400 gamma=32'd1;row=32'd227;
#400 gamma=32'd1;row=32'd123;
#400 gamma=32'd4;row=32'd419;
#400 gamma=32'd3;row=32'd120;
#400 gamma=32'd1;row=32'd274;
#400 gamma=32'd5;row=32'd403;
#400 gamma=32'd5;row=32'd126;
#400 gamma=32'd2;row=32'd243;
#400 gamma=32'd1;row=32'd242;
#400 gamma=32'd3;row=32'd210;
#400 gamma=32'd5;row=32'd548;
#400 gamma=32'd2;row=32'd537;
#400 gamma=32'd2;row=32'd340;
#400 gamma=32'd1;row=32'd359;
#400 gamma=32'd5;row=32'd555;
#400 gamma=32'd2;row=32'd141;
#400 gamma=32'd4;row=32'd92;
#400 gamma=32'd5;row=32'd285;
#400 gamma=32'd3;row=32'd498;
#400 gamma=32'd4;row=32'd21;
#400 gamma=32'd4;row=32'd445;
#400 gamma=32'd5;row=32'd399;
#400 gamma=32'd2;row=32'd124;
#400 gamma=32'd1;row=32'd305;
#400 gamma=32'd3;row=32'd308;
#400 gamma=32'd3;row=32'd276;
#400 gamma=32'd2;row=32'd6;
#400 gamma=32'd5;row=32'd397;
#400 gamma=32'd1;row=32'd426;
#400 gamma=32'd3;row=32'd410;
#400 gamma=32'd1;row=32'd238;
#400 gamma=32'd4;row=32'd328;
#400 gamma=32'd3;row=32'd103;
#400 gamma=32'd2;row=32'd447;
#400 gamma=32'd2;row=32'd398;
#400 gamma=32'd4;row=32'd31;
#400 gamma=32'd4;row=32'd464;
#400 gamma=32'd3;row=32'd293;
#400 gamma=32'd2;row=32'd385;
#400 gamma=32'd4;row=32'd94;
#400 gamma=32'd5;row=32'd473;
#400 gamma=32'd5;row=32'd373;
#400 gamma=32'd5;row=32'd435;
#400 gamma=32'd3;row=32'd507;
#400 gamma=32'd1;row=32'd374;
#400 gamma=32'd5;row=32'd442;
#400 gamma=32'd2;row=32'd451;
#400 gamma=32'd5;row=32'd274;
#400 gamma=32'd4;row=32'd9;
#400 gamma=32'd3;row=32'd182;
#400 gamma=32'd3;row=32'd365;
#400 gamma=32'd1;row=32'd172;
#400 gamma=32'd5;row=32'd119;
#400 gamma=32'd4;row=32'd299;
#400 gamma=32'd4;row=32'd505;
#400 gamma=32'd5;row=32'd51;
#400 gamma=32'd3;row=32'd262;
#400 gamma=32'd4;row=32'd151;
#400 gamma=32'd5;row=32'd511;
#400 gamma=32'd1;row=32'd327;
#400 gamma=32'd1;row=32'd240;
#400 gamma=32'd4;row=32'd159;
#400 gamma=32'd2;row=32'd38;
#400 gamma=32'd5;row=32'd527;
#400 gamma=32'd1;row=32'd343;
#400 gamma=32'd3;row=32'd347;
#400 gamma=32'd5;row=32'd493;
#400 gamma=32'd2;row=32'd363;
#400 gamma=32'd3;row=32'd536;
#400 gamma=32'd1;row=32'd515;
#400 gamma=32'd4;row=32'd415;
#400 gamma=32'd1;row=32'd45;
#400 gamma=32'd2;row=32'd118;
#400 gamma=32'd4;row=32'd248;
#400 gamma=32'd3;row=32'd284;
#400 gamma=32'd5;row=32'd234;
#400 gamma=32'd5;row=32'd330;
#400 gamma=32'd4;row=32'd294;
#400 gamma=32'd5;row=32'd154;
#400 gamma=32'd1;row=32'd266;
#400 gamma=32'd4;row=32'd235;
#400 gamma=32'd4;row=32'd432;
#400 gamma=32'd1;row=32'd39;
#400 gamma=32'd4;row=32'd119;
#400 gamma=32'd2;row=32'd520;
#400 gamma=32'd3;row=32'd311;
#400 gamma=32'd4;row=32'd293;
#400 gamma=32'd4;row=32'd506;
#400 gamma=32'd1;row=32'd308;
#400 gamma=32'd2;row=32'd3;
#400 gamma=32'd5;row=32'd72;
#400 gamma=32'd4;row=32'd224;
#400 gamma=32'd4;row=32'd551;
#400 gamma=32'd1;row=32'd486;
#400 gamma=32'd1;row=32'd449;
#400 gamma=32'd4;row=32'd179;
#400 gamma=32'd4;row=32'd263;
#400 gamma=32'd4;row=32'd15;
#400 gamma=32'd4;row=32'd87;
#400 gamma=32'd3;row=32'd224;
#400 gamma=32'd3;row=32'd262;
#400 gamma=32'd4;row=32'd89;
#400 gamma=32'd4;row=32'd333;
#400 gamma=32'd2;row=32'd460;
#400 gamma=32'd2;row=32'd401;
#400 gamma=32'd5;row=32'd310;
#400 gamma=32'd4;row=32'd464;
#400 gamma=32'd5;row=32'd141;
#400 gamma=32'd3;row=32'd489;
#400 gamma=32'd4;row=32'd128;
#400 gamma=32'd2;row=32'd461;
#400 gamma=32'd3;row=32'd65;
#400 gamma=32'd3;row=32'd163;
#400 gamma=32'd2;row=32'd335;
#400 gamma=32'd3;row=32'd75;
#400 gamma=32'd5;row=32'd482;
#400 gamma=32'd3;row=32'd290;
#400 gamma=32'd2;row=32'd448;
#400 gamma=32'd3;row=32'd230;
#400 gamma=32'd2;row=32'd294;
#400 gamma=32'd2;row=32'd393;
#400 gamma=32'd1;row=32'd457;
#400 gamma=32'd2;row=32'd489;
#400 gamma=32'd5;row=32'd330;
#400 gamma=32'd5;row=32'd393;
#400 gamma=32'd1;row=32'd447;
#400 gamma=32'd1;row=32'd124;
#400 gamma=32'd2;row=32'd6;
#400 gamma=32'd2;row=32'd157;
#400 gamma=32'd5;row=32'd187;
#400 gamma=32'd1;row=32'd379;
#400 gamma=32'd3;row=32'd129;
#400 gamma=32'd2;row=32'd75;
#400 gamma=32'd2;row=32'd520;
#400 gamma=32'd5;row=32'd241;
#400 gamma=32'd1;row=32'd550;
#400 gamma=32'd1;row=32'd534;
#400 gamma=32'd1;row=32'd484;
#400 gamma=32'd4;row=32'd16;
#400 gamma=32'd3;row=32'd132;
#400 gamma=32'd5;row=32'd222;
#400 gamma=32'd4;row=32'd522;
#400 gamma=32'd4;row=32'd534;
#400 gamma=32'd3;row=32'd516;
#400 gamma=32'd1;row=32'd57;
#400 gamma=32'd5;row=32'd38;
#400 gamma=32'd5;row=32'd149;
#400 gamma=32'd2;row=32'd496;
#400 gamma=32'd5;row=32'd287;
#400 gamma=32'd2;row=32'd315;
#400 gamma=32'd2;row=32'd460;
#400 gamma=32'd4;row=32'd191;
#400 gamma=32'd5;row=32'd218;
#400 gamma=32'd3;row=32'd14;
#400 gamma=32'd4;row=32'd256;
#400 gamma=32'd5;row=32'd6;
#400 gamma=32'd4;row=32'd32;
#400 gamma=32'd5;row=32'd182;
#400 gamma=32'd3;row=32'd465;
#400 gamma=32'd1;row=32'd273;
#400 gamma=32'd3;row=32'd139;
#400 gamma=32'd5;row=32'd58;
#400 gamma=32'd4;row=32'd369;
#400 gamma=32'd2;row=32'd519;
#400 gamma=32'd5;row=32'd442;
#400 gamma=32'd2;row=32'd525;
#400 gamma=32'd4;row=32'd88;
#400 gamma=32'd1;row=32'd243;
#400 gamma=32'd4;row=32'd40;
#400 gamma=32'd3;row=32'd267;
#400 gamma=32'd4;row=32'd430;
#400 gamma=32'd4;row=32'd396;
#400 gamma=32'd3;row=32'd182;
#400 gamma=32'd5;row=32'd27;
#400 gamma=32'd1;row=32'd83;
#400 gamma=32'd2;row=32'd354;
#400 gamma=32'd3;row=32'd256;
#400 gamma=32'd3;row=32'd159;
#400 gamma=32'd2;row=32'd428;
#400 gamma=32'd2;row=32'd124;
#400 gamma=32'd3;row=32'd177;
#400 gamma=32'd4;row=32'd450;
#400 gamma=32'd4;row=32'd323;
#400 gamma=32'd2;row=32'd73;
#400 gamma=32'd2;row=32'd544;
#400 gamma=32'd3;row=32'd464;
#400 gamma=32'd4;row=32'd430;
#400 gamma=32'd2;row=32'd224;
#400 gamma=32'd2;row=32'd164;
#400 gamma=32'd5;row=32'd458;
#400 gamma=32'd2;row=32'd449;
#400 gamma=32'd1;row=32'd80;
#400 gamma=32'd3;row=32'd545;
#400 gamma=32'd3;row=32'd25;
#400 gamma=32'd2;row=32'd248;
#400 gamma=32'd5;row=32'd176;
#400 gamma=32'd4;row=32'd522;
#400 gamma=32'd5;row=32'd155;
#400 gamma=32'd3;row=32'd220;
#400 gamma=32'd2;row=32'd173;
#400 gamma=32'd4;row=32'd335;
#400 gamma=32'd1;row=32'd555;
#400 gamma=32'd1;row=32'd87;
#400 gamma=32'd4;row=32'd401;
#400 gamma=32'd1;row=32'd201;
#400 gamma=32'd2;row=32'd410;
#400 gamma=32'd5;row=32'd265;
#400 gamma=32'd4;row=32'd334;
#400 gamma=32'd2;row=32'd305;
#400 gamma=32'd3;row=32'd240;
#400 gamma=32'd4;row=32'd34;
#400 gamma=32'd4;row=32'd227;
#400 gamma=32'd5;row=32'd40;
#400 gamma=32'd4;row=32'd263;
#400 gamma=32'd2;row=32'd477;
#400 gamma=32'd2;row=32'd344;
#400 gamma=32'd1;row=32'd403;
#400 gamma=32'd4;row=32'd287;
#400 gamma=32'd5;row=32'd453;
#400 gamma=32'd5;row=32'd29;
#400 gamma=32'd4;row=32'd207;
#400 gamma=32'd3;row=32'd181;
#400 gamma=32'd2;row=32'd521;
#400 gamma=32'd2;row=32'd103;
#400 gamma=32'd4;row=32'd59;
#400 gamma=32'd1;row=32'd296;
#400 gamma=32'd2;row=32'd322;
#400 gamma=32'd1;row=32'd29;
#400 gamma=32'd2;row=32'd434;
#400 gamma=32'd2;row=32'd513;
#400 gamma=32'd3;row=32'd121;
#400 gamma=32'd2;row=32'd129;
#400 gamma=32'd4;row=32'd413;
#400 gamma=32'd2;row=32'd260;
#400 gamma=32'd2;row=32'd67;
#400 gamma=32'd3;row=32'd365;
#400 gamma=32'd4;row=32'd397;
#400 gamma=32'd2;row=32'd409;
#400 gamma=32'd5;row=32'd492;
#400 gamma=32'd1;row=32'd102;
#400 gamma=32'd3;row=32'd84;
#400 gamma=32'd1;row=32'd103;
#400 gamma=32'd3;row=32'd526;
#400 gamma=32'd4;row=32'd137;
#400 gamma=32'd3;row=32'd189;
#400 gamma=32'd1;row=32'd2;
#400 gamma=32'd2;row=32'd489;
#400 gamma=32'd4;row=32'd174;
#400 gamma=32'd1;row=32'd179;
#400 gamma=32'd3;row=32'd55;
#400 gamma=32'd3;row=32'd311;
#400 gamma=32'd2;row=32'd337;
#400 gamma=32'd1;row=32'd89;
#400 gamma=32'd3;row=32'd286;
#400 gamma=32'd4;row=32'd439;
#400 gamma=32'd5;row=32'd559;
#400 gamma=32'd3;row=32'd513;
#400 gamma=32'd5;row=32'd518;
#400 gamma=32'd3;row=32'd187;
#400 gamma=32'd1;row=32'd271;
#400 gamma=32'd1;row=32'd319;
#400 gamma=32'd1;row=32'd421;
#400 gamma=32'd1;row=32'd439;
#400 gamma=32'd4;row=32'd519;
#400 gamma=32'd2;row=32'd93;
#400 gamma=32'd1;row=32'd44;
#400 gamma=32'd4;row=32'd249;
#400 gamma=32'd2;row=32'd524;
#400 gamma=32'd2;row=32'd304;
#400 gamma=32'd3;row=32'd400;
#400 gamma=32'd2;row=32'd33;
#400 gamma=32'd3;row=32'd260;
#400 gamma=32'd2;row=32'd192;
#400 gamma=32'd2;row=32'd427;
#400 gamma=32'd1;row=32'd454;
#400 gamma=32'd3;row=32'd501;
#400 gamma=32'd3;row=32'd198;
#400 gamma=32'd3;row=32'd27;
#400 gamma=32'd2;row=32'd263;
#400 gamma=32'd5;row=32'd310;
#400 gamma=32'd5;row=32'd37;
#400 gamma=32'd1;row=32'd454;
#400 gamma=32'd3;row=32'd389;
#400 gamma=32'd3;row=32'd165;
#400 gamma=32'd3;row=32'd94;
#400 gamma=32'd4;row=32'd392;
#400 gamma=32'd5;row=32'd158;
#400 gamma=32'd3;row=32'd497;
#400 gamma=32'd2;row=32'd190;
#400 gamma=32'd1;row=32'd494;
#400 gamma=32'd2;row=32'd518;
#400 gamma=32'd4;row=32'd427;
#400 gamma=32'd2;row=32'd542;
#400 gamma=32'd4;row=32'd373;
#400 gamma=32'd1;row=32'd479;
#400 gamma=32'd5;row=32'd412;
#400 gamma=32'd5;row=32'd179;
#400 gamma=32'd5;row=32'd499;
#400 gamma=32'd3;row=32'd535;
#400 gamma=32'd5;row=32'd555;
#400 gamma=32'd1;row=32'd210;
#400 gamma=32'd2;row=32'd384;
#400 gamma=32'd2;row=32'd559;
#400 gamma=32'd4;row=32'd377;
#400 gamma=32'd2;row=32'd33;
#400 gamma=32'd4;row=32'd255;
#400 gamma=32'd2;row=32'd364;
#400 gamma=32'd4;row=32'd26;
#400 gamma=32'd3;row=32'd205;
#400 gamma=32'd2;row=32'd218;
#400 gamma=32'd1;row=32'd170;
#400 gamma=32'd3;row=32'd33;
#400 gamma=32'd4;row=32'd538;
#400 gamma=32'd1;row=32'd375;
#400 gamma=32'd2;row=32'd37;
#400 gamma=32'd1;row=32'd342;
#400 gamma=32'd1;row=32'd143;
#400 gamma=32'd5;row=32'd415;
#400 gamma=32'd4;row=32'd344;
#400 gamma=32'd4;row=32'd370;
#400 gamma=32'd4;row=32'd62;
#400 gamma=32'd5;row=32'd223;
#400 gamma=32'd4;row=32'd2;
#400 gamma=32'd1;row=32'd363;
#400 gamma=32'd5;row=32'd431;
#400 gamma=32'd2;row=32'd158;
#400 gamma=32'd4;row=32'd269;
#400 gamma=32'd3;row=32'd172;
#400 gamma=32'd5;row=32'd87;
#400 gamma=32'd1;row=32'd350;
#400 gamma=32'd3;row=32'd445;
#400 gamma=32'd4;row=32'd383;
#400 gamma=32'd5;row=32'd346;
#400 gamma=32'd4;row=32'd473;
#400 gamma=32'd5;row=32'd370;
#400 gamma=32'd3;row=32'd348;
#400 gamma=32'd5;row=32'd215;
#400 gamma=32'd2;row=32'd302;
#400 gamma=32'd2;row=32'd315;
#400 gamma=32'd5;row=32'd129;
#400 gamma=32'd2;row=32'd452;
#400 gamma=32'd1;row=32'd394;
#400 gamma=32'd3;row=32'd459;
#400 gamma=32'd2;row=32'd27;
#400 gamma=32'd5;row=32'd155;
#400 gamma=32'd3;row=32'd56;
#400 gamma=32'd4;row=32'd366;
#400 gamma=32'd1;row=32'd129;
#400 gamma=32'd2;row=32'd69;
#400 gamma=32'd4;row=32'd509;
#400 gamma=32'd5;row=32'd327;
#400 gamma=32'd5;row=32'd291;
#400 gamma=32'd3;row=32'd137;
#400 gamma=32'd1;row=32'd412;
#400 gamma=32'd4;row=32'd292;
#400 gamma=32'd1;row=32'd419;
#400 gamma=32'd5;row=32'd287;
#400 gamma=32'd1;row=32'd505;
#400 gamma=32'd1;row=32'd550;
#400 gamma=32'd2;row=32'd307;
#400 gamma=32'd2;row=32'd444;
#400 gamma=32'd5;row=32'd300;
#400 gamma=32'd3;row=32'd268;
#400 gamma=32'd2;row=32'd132;
#400 gamma=32'd3;row=32'd129;
#400 gamma=32'd5;row=32'd74;
#400 gamma=32'd4;row=32'd529;
#400 gamma=32'd4;row=32'd180;
#400 gamma=32'd1;row=32'd499;
#400 gamma=32'd2;row=32'd462;
#400 gamma=32'd4;row=32'd332;
#400 gamma=32'd2;row=32'd485;
#400 gamma=32'd5;row=32'd176;
#400 gamma=32'd4;row=32'd357;
#400 gamma=32'd3;row=32'd491;
#400 gamma=32'd2;row=32'd203;
#400 gamma=32'd3;row=32'd23;
#400 gamma=32'd2;row=32'd38;
#400 gamma=32'd1;row=32'd175;
#400 gamma=32'd2;row=32'd547;
#400 gamma=32'd4;row=32'd505;
#400 gamma=32'd3;row=32'd4;
#400 gamma=32'd3;row=32'd121;
#400 gamma=32'd3;row=32'd341;
#400 gamma=32'd5;row=32'd343;
#400 gamma=32'd1;row=32'd519;
#400 gamma=32'd4;row=32'd510;
#400 gamma=32'd4;row=32'd3;
#400 gamma=32'd3;row=32'd200;
#400 gamma=32'd4;row=32'd340;
#400 gamma=32'd4;row=32'd0;
#400 gamma=32'd3;row=32'd212;
#400 gamma=32'd3;row=32'd153;
#400 gamma=32'd3;row=32'd102;
#400 gamma=32'd4;row=32'd365;
#400 gamma=32'd5;row=32'd408;
#400 gamma=32'd5;row=32'd236;
#400 gamma=32'd1;row=32'd430;
#400 gamma=32'd1;row=32'd271;
#400 gamma=32'd2;row=32'd517;
#400 gamma=32'd3;row=32'd37;
#400 gamma=32'd4;row=32'd325;
#400 gamma=32'd3;row=32'd322;
#400 gamma=32'd2;row=32'd74;
#400 gamma=32'd4;row=32'd487;
#400 gamma=32'd3;row=32'd479;
#400 gamma=32'd3;row=32'd97;
#400 gamma=32'd2;row=32'd378;
#400 gamma=32'd3;row=32'd101;
#400 gamma=32'd3;row=32'd494;
#400 gamma=32'd3;row=32'd69;
#400 gamma=32'd3;row=32'd105;
#400 gamma=32'd3;row=32'd466;
#400 gamma=32'd4;row=32'd327;
#400 gamma=32'd5;row=32'd364;
#400 gamma=32'd5;row=32'd167;
#400 gamma=32'd1;row=32'd367;
#400 gamma=32'd4;row=32'd495;
#400 gamma=32'd3;row=32'd482;
#400 gamma=32'd2;row=32'd479;
#400 gamma=32'd2;row=32'd126;
#400 gamma=32'd4;row=32'd92;
#400 gamma=32'd3;row=32'd547;
#400 gamma=32'd2;row=32'd510;
#400 gamma=32'd5;row=32'd374;
#400 gamma=32'd2;row=32'd450;
#400 gamma=32'd4;row=32'd170;
#400 gamma=32'd2;row=32'd130;
#400 gamma=32'd5;row=32'd224;
#400 gamma=32'd2;row=32'd287;
#400 gamma=32'd3;row=32'd81;
#400 gamma=32'd2;row=32'd313;
#400 gamma=32'd2;row=32'd552;
#400 gamma=32'd2;row=32'd102;
#400 gamma=32'd5;row=32'd308;
#400 gamma=32'd1;row=32'd514;
#400 gamma=32'd2;row=32'd318;
#400 gamma=32'd3;row=32'd187;
#400 gamma=32'd1;row=32'd127;
#400 gamma=32'd4;row=32'd170;
#400 gamma=32'd3;row=32'd228;
#400 gamma=32'd3;row=32'd223;
#400 gamma=32'd2;row=32'd354;
#400 gamma=32'd2;row=32'd40;
#400 gamma=32'd2;row=32'd212;
#400 gamma=32'd2;row=32'd400;
#400 gamma=32'd2;row=32'd441;
#400 gamma=32'd1;row=32'd417;
#400 gamma=32'd2;row=32'd400;
#400 gamma=32'd5;row=32'd160;
#400 gamma=32'd1;row=32'd328;
#400 gamma=32'd2;row=32'd146;
#400 gamma=32'd5;row=32'd557;
#400 gamma=32'd4;row=32'd93;
#400 gamma=32'd4;row=32'd100;
#400 gamma=32'd3;row=32'd113;
#400 gamma=32'd2;row=32'd495;
#400 gamma=32'd3;row=32'd233;
#400 gamma=32'd4;row=32'd67;
#400 gamma=32'd1;row=32'd249;
#400 gamma=32'd3;row=32'd449;
#400 gamma=32'd1;row=32'd372;
#400 gamma=32'd3;row=32'd468;
#400 gamma=32'd4;row=32'd319;
#400 gamma=32'd5;row=32'd166;
#400 gamma=32'd5;row=32'd478;
#400 gamma=32'd1;row=32'd242;
#400 gamma=32'd4;row=32'd447;
#400 gamma=32'd4;row=32'd500;
#400 gamma=32'd4;row=32'd499;
#400 gamma=32'd4;row=32'd153;
#400 gamma=32'd5;row=32'd531;
#400 gamma=32'd2;row=32'd76;
#400 gamma=32'd2;row=32'd235;
#400 gamma=32'd2;row=32'd386;
#400 gamma=32'd4;row=32'd112;
#400 gamma=32'd1;row=32'd406;
#400 gamma=32'd3;row=32'd308;
#400 gamma=32'd3;row=32'd262;
#400 gamma=32'd4;row=32'd427;
#400 gamma=32'd5;row=32'd527;
#400 gamma=32'd2;row=32'd340;
#400 gamma=32'd5;row=32'd265;
#400 gamma=32'd1;row=32'd208;
#400 gamma=32'd4;row=32'd327;
#400 gamma=32'd3;row=32'd187;
#400 gamma=32'd1;row=32'd527;
#400 gamma=32'd5;row=32'd510;
#400 gamma=32'd2;row=32'd333;
#400 gamma=32'd4;row=32'd457;
#400 gamma=32'd1;row=32'd110;
#400 gamma=32'd5;row=32'd166;
#400 gamma=32'd2;row=32'd165;
#400 gamma=32'd5;row=32'd274;
#400 gamma=32'd2;row=32'd218;
#400 gamma=32'd3;row=32'd170;
#400 gamma=32'd5;row=32'd114;
#400 gamma=32'd1;row=32'd542;
#400 gamma=32'd1;row=32'd104;
#400 gamma=32'd2;row=32'd72;
#400 gamma=32'd5;row=32'd438;
#400 gamma=32'd3;row=32'd128;
#400 gamma=32'd4;row=32'd320;
#400 gamma=32'd5;row=32'd432;
#400 gamma=32'd4;row=32'd80;
#400 gamma=32'd3;row=32'd210;
#400 gamma=32'd2;row=32'd528;
#400 gamma=32'd3;row=32'd128;
#400 gamma=32'd1;row=32'd192;
#400 gamma=32'd3;row=32'd251;
#400 gamma=32'd1;row=32'd247;
#400 gamma=32'd4;row=32'd385;
#400 gamma=32'd5;row=32'd45;
#400 gamma=32'd3;row=32'd83;
#400 gamma=32'd2;row=32'd544;
#400 gamma=32'd5;row=32'd464;
#400 gamma=32'd1;row=32'd482;
#400 gamma=32'd1;row=32'd13;
#400 gamma=32'd3;row=32'd213;
#400 gamma=32'd4;row=32'd505;
#400 gamma=32'd5;row=32'd453;
#400 gamma=32'd2;row=32'd302;
#400 gamma=32'd1;row=32'd86;
#400 gamma=32'd3;row=32'd425;
#400 gamma=32'd4;row=32'd224;
#400 gamma=32'd3;row=32'd123;
#400 gamma=32'd1;row=32'd524;
#400 gamma=32'd3;row=32'd511;
#400 gamma=32'd2;row=32'd358;
#400 gamma=32'd5;row=32'd357;
#400 gamma=32'd1;row=32'd111;
#400 gamma=32'd4;row=32'd374;
#400 gamma=32'd3;row=32'd255;
#400 gamma=32'd3;row=32'd248;
#400 gamma=32'd2;row=32'd415;
#400 gamma=32'd3;row=32'd98;
#400 gamma=32'd3;row=32'd142;
#400 gamma=32'd2;row=32'd250;
#400 gamma=32'd2;row=32'd88;
#400 gamma=32'd3;row=32'd314;
#400 gamma=32'd5;row=32'd427;
#400 gamma=32'd2;row=32'd536;
#400 gamma=32'd4;row=32'd468;
#400 gamma=32'd5;row=32'd153;
#400 gamma=32'd5;row=32'd7;
#400 gamma=32'd3;row=32'd286;
#400 gamma=32'd4;row=32'd450;
#400 gamma=32'd4;row=32'd306;
#400 gamma=32'd2;row=32'd470;
#400 gamma=32'd2;row=32'd222;
#400 gamma=32'd3;row=32'd438;
#400 gamma=32'd1;row=32'd472;
#400 gamma=32'd2;row=32'd507;
#400 gamma=32'd3;row=32'd89;
#400 gamma=32'd1;row=32'd349;
#400 gamma=32'd3;row=32'd18;
#400 gamma=32'd4;row=32'd78;
#400 gamma=32'd5;row=32'd243;
#400 gamma=32'd1;row=32'd76;
#400 gamma=32'd4;row=32'd156;
#400 gamma=32'd2;row=32'd65;
#400 gamma=32'd1;row=32'd37;
#400 gamma=32'd5;row=32'd480;
#400 gamma=32'd4;row=32'd180;
#400 gamma=32'd4;row=32'd446;
#400 gamma=32'd2;row=32'd401;
#400 gamma=32'd1;row=32'd417;
#400 gamma=32'd1;row=32'd169;
#400 gamma=32'd5;row=32'd208;
#400 gamma=32'd5;row=32'd1;
#400 gamma=32'd4;row=32'd108;
#400 gamma=32'd2;row=32'd250;
#400 gamma=32'd5;row=32'd276;
#400 gamma=32'd5;row=32'd558;
#400 gamma=32'd2;row=32'd399;
#400 gamma=32'd4;row=32'd428;
#400 gamma=32'd3;row=32'd149;
#400 gamma=32'd5;row=32'd325;
#400 gamma=32'd5;row=32'd248;
#400 gamma=32'd3;row=32'd254;
#400 gamma=32'd1;row=32'd381;
#400 gamma=32'd1;row=32'd402;
#400 gamma=32'd5;row=32'd325;
#400 gamma=32'd1;row=32'd451;
#400 gamma=32'd1;row=32'd456;
#400 gamma=32'd1;row=32'd313;
#400 gamma=32'd4;row=32'd249;
#400 gamma=32'd3;row=32'd152;
#400 gamma=32'd4;row=32'd426;
#400 gamma=32'd3;row=32'd425;
#400 gamma=32'd3;row=32'd548;
#400 gamma=32'd5;row=32'd76;
#400 gamma=32'd2;row=32'd169;
#400 gamma=32'd1;row=32'd229;
#400 gamma=32'd2;row=32'd230;
#400 gamma=32'd3;row=32'd559;
#400 gamma=32'd1;row=32'd277;
#400 gamma=32'd5;row=32'd28;
#400 gamma=32'd4;row=32'd157;
#400 gamma=32'd3;row=32'd287;
#400 gamma=32'd5;row=32'd263;
#400 gamma=32'd3;row=32'd200;
#400 gamma=32'd1;row=32'd418;
#400 gamma=32'd5;row=32'd342;
#400 gamma=32'd1;row=32'd443;
#400 gamma=32'd2;row=32'd316;
#400 gamma=32'd3;row=32'd494;
#400 gamma=32'd4;row=32'd532;
#400 gamma=32'd3;row=32'd124;
#400 gamma=32'd4;row=32'd205;
#400 gamma=32'd3;row=32'd10;
#400 gamma=32'd4;row=32'd248;
#400 gamma=32'd5;row=32'd476;
#400 gamma=32'd1;row=32'd4;
#400 gamma=32'd4;row=32'd247;
#400 gamma=32'd3;row=32'd37;
#400 gamma=32'd3;row=32'd305;
#400 gamma=32'd4;row=32'd511;
#400 gamma=32'd2;row=32'd243;
#400 gamma=32'd2;row=32'd24;
#400 gamma=32'd5;row=32'd541;
#400 gamma=32'd1;row=32'd181;
#400 gamma=32'd3;row=32'd246;
#400 gamma=32'd4;row=32'd192;
#400 gamma=32'd5;row=32'd58;
#400 gamma=32'd5;row=32'd92;
#400 gamma=32'd4;row=32'd41;
#400 gamma=32'd3;row=32'd143;
#400 gamma=32'd2;row=32'd374;
#400 gamma=32'd3;row=32'd85;
#400 gamma=32'd5;row=32'd180;
#400 gamma=32'd2;row=32'd36;
#400 gamma=32'd1;row=32'd393;
#400 gamma=32'd5;row=32'd208;
#400 gamma=32'd1;row=32'd262;
#400 gamma=32'd1;row=32'd62;
#400 gamma=32'd4;row=32'd399;
#400 gamma=32'd4;row=32'd212;
#400 gamma=32'd3;row=32'd66;
#400 gamma=32'd2;row=32'd481;
#400 gamma=32'd1;row=32'd133;
#400 gamma=32'd3;row=32'd235;
#400 gamma=32'd1;row=32'd433;
#400 gamma=32'd5;row=32'd183;
#400 gamma=32'd5;row=32'd507;
#400 gamma=32'd5;row=32'd311;
#400 gamma=32'd4;row=32'd195;
#400 gamma=32'd4;row=32'd339;
#400 gamma=32'd4;row=32'd151;
#400 gamma=32'd3;row=32'd51;
#400 gamma=32'd3;row=32'd460;
#400 gamma=32'd4;row=32'd51;
#400 gamma=32'd5;row=32'd438;
#400 gamma=32'd4;row=32'd9;
#400 gamma=32'd5;row=32'd390;
#400 gamma=32'd1;row=32'd206;
#400 gamma=32'd3;row=32'd129;
#400 gamma=32'd1;row=32'd170;
#400 gamma=32'd3;row=32'd512;
#400 gamma=32'd1;row=32'd173;
#400 gamma=32'd5;row=32'd511;
#400 gamma=32'd1;row=32'd275;
#400 gamma=32'd5;row=32'd115;
#400 gamma=32'd3;row=32'd296;
#400 gamma=32'd3;row=32'd108;
#400 gamma=32'd3;row=32'd435;
#400 gamma=32'd3;row=32'd166;
#400 gamma=32'd4;row=32'd321;
#400 gamma=32'd4;row=32'd350;
#400 gamma=32'd1;row=32'd281;
#400 gamma=32'd4;row=32'd112;
#400 gamma=32'd2;row=32'd39;
#400 gamma=32'd1;row=32'd262;
#400 gamma=32'd3;row=32'd8;
#400 gamma=32'd5;row=32'd188;
#400 gamma=32'd4;row=32'd440;
#400 gamma=32'd5;row=32'd315;
#400 gamma=32'd2;row=32'd395;
#400 gamma=32'd3;row=32'd367;
#400 gamma=32'd5;row=32'd377;
#400 gamma=32'd4;row=32'd514;
#400 gamma=32'd4;row=32'd547;
#400 gamma=32'd2;row=32'd262;
#400 gamma=32'd5;row=32'd292;
#400 gamma=32'd4;row=32'd223;
#400 gamma=32'd5;row=32'd67;
#400 gamma=32'd5;row=32'd71;
#400 gamma=32'd5;row=32'd335;
#400 gamma=32'd2;row=32'd495;
#400 gamma=32'd4;row=32'd323;
#400 gamma=32'd2;row=32'd87;
#400 gamma=32'd4;row=32'd236;
#400 gamma=32'd4;row=32'd390;
#400 gamma=32'd3;row=32'd258;
#400 gamma=32'd5;row=32'd0;
#400 gamma=32'd4;row=32'd186;
#400 gamma=32'd1;row=32'd58;
#400 gamma=32'd2;row=32'd448;
#400 gamma=32'd4;row=32'd306;
#400 gamma=32'd3;row=32'd233;
#400 gamma=32'd1;row=32'd493;
#400 gamma=32'd4;row=32'd390;
#400 gamma=32'd3;row=32'd443;
#400 gamma=32'd2;row=32'd104;
#400 gamma=32'd3;row=32'd538;
#400 gamma=32'd1;row=32'd86;
#400 gamma=32'd2;row=32'd38;
#400 gamma=32'd4;row=32'd138;
#400 gamma=32'd4;row=32'd30;
#400 gamma=32'd3;row=32'd448;
#400 gamma=32'd2;row=32'd382;
#400 gamma=32'd3;row=32'd385;
#400 gamma=32'd5;row=32'd266;
#400 gamma=32'd1;row=32'd277;
#400 gamma=32'd2;row=32'd330;
#400 gamma=32'd3;row=32'd363;
#400 gamma=32'd5;row=32'd162;
#400 gamma=32'd1;row=32'd532;
#400 gamma=32'd5;row=32'd196;
#400 gamma=32'd5;row=32'd529;
#400 gamma=32'd5;row=32'd184;
#400 gamma=32'd4;row=32'd92;
#400 gamma=32'd3;row=32'd486;
#400 gamma=32'd2;row=32'd176;
#400 gamma=32'd2;row=32'd276;
#400 gamma=32'd4;row=32'd265;
#400 gamma=32'd2;row=32'd512;
#400 gamma=32'd5;row=32'd392;
#400 gamma=32'd1;row=32'd345;
#400 gamma=32'd4;row=32'd186;
#400 gamma=32'd5;row=32'd138;
#400 gamma=32'd5;row=32'd34;
#400 gamma=32'd1;row=32'd268;
#400 gamma=32'd3;row=32'd452;
#400 gamma=32'd5;row=32'd242;
#400 gamma=32'd4;row=32'd518;
#400 gamma=32'd3;row=32'd94;
#400 gamma=32'd4;row=32'd189;
#400 gamma=32'd1;row=32'd44;
#400 gamma=32'd1;row=32'd541;
#400 gamma=32'd2;row=32'd50;
#400 gamma=32'd3;row=32'd377;
#400 gamma=32'd3;row=32'd479;
#400 gamma=32'd5;row=32'd430;
#400 gamma=32'd5;row=32'd147;
#400 gamma=32'd4;row=32'd392;
#400 gamma=32'd5;row=32'd26;
#400 gamma=32'd3;row=32'd381;
#400 gamma=32'd2;row=32'd0;
#400 gamma=32'd1;row=32'd540;
#400 gamma=32'd5;row=32'd445;
#400 gamma=32'd4;row=32'd440;
#400 gamma=32'd5;row=32'd48;
#400 gamma=32'd2;row=32'd512;
#400 gamma=32'd4;row=32'd419;
#400 gamma=32'd1;row=32'd258;
#400 gamma=32'd3;row=32'd460;
#400 gamma=32'd5;row=32'd333;
#400 gamma=32'd1;row=32'd499;
#400 gamma=32'd5;row=32'd58;
#400 gamma=32'd2;row=32'd297;
#400 gamma=32'd3;row=32'd116;
#400 gamma=32'd1;row=32'd240;
#400 gamma=32'd4;row=32'd149;
#400 gamma=32'd1;row=32'd443;
#400 gamma=32'd4;row=32'd536;
#400 gamma=32'd3;row=32'd364;
#400 gamma=32'd4;row=32'd527;
#400 gamma=32'd3;row=32'd425;
#400 gamma=32'd5;row=32'd393;
#400 gamma=32'd1;row=32'd153;
#400 gamma=32'd1;row=32'd413;
#400 gamma=32'd1;row=32'd416;
#400 gamma=32'd1;row=32'd9;
#400 gamma=32'd1;row=32'd381;
#400 gamma=32'd3;row=32'd354;
#400 gamma=32'd1;row=32'd322;
#400 gamma=32'd5;row=32'd121;
#400 gamma=32'd3;row=32'd499;
#400 gamma=32'd5;row=32'd379;
#400 gamma=32'd3;row=32'd340;
#400 gamma=32'd3;row=32'd444;
#400 gamma=32'd2;row=32'd170;
#400 gamma=32'd3;row=32'd68;
#400 gamma=32'd1;row=32'd284;
#400 gamma=32'd2;row=32'd44;
#400 gamma=32'd1;row=32'd89;
#400 gamma=32'd3;row=32'd346;
#400 gamma=32'd1;row=32'd379;
#400 gamma=32'd2;row=32'd443;
#400 gamma=32'd1;row=32'd473;
#400 gamma=32'd4;row=32'd503;
#400 gamma=32'd5;row=32'd465;
#400 gamma=32'd1;row=32'd200;
#400 gamma=32'd5;row=32'd73;
#400 gamma=32'd3;row=32'd165;
#400 gamma=32'd2;row=32'd286;
#400 gamma=32'd5;row=32'd7;
#400 gamma=32'd2;row=32'd144;
#400 gamma=32'd5;row=32'd415;
#400 gamma=32'd1;row=32'd225;
#400 gamma=32'd5;row=32'd111;
#400 gamma=32'd2;row=32'd7;
#400 gamma=32'd1;row=32'd331;
#400 gamma=32'd4;row=32'd17;
#400 gamma=32'd4;row=32'd279;
#400 gamma=32'd2;row=32'd111;
#400 gamma=32'd5;row=32'd64;
#400 gamma=32'd4;row=32'd288;
#400 gamma=32'd3;row=32'd8;
#400 gamma=32'd4;row=32'd77;
#400 gamma=32'd3;row=32'd389;
#400 gamma=32'd2;row=32'd89;
#400 gamma=32'd2;row=32'd176;
#400 gamma=32'd5;row=32'd101;
#400 gamma=32'd3;row=32'd15;
#400 gamma=32'd2;row=32'd146;
#400 gamma=32'd2;row=32'd400;
#400 gamma=32'd3;row=32'd246;
#400 gamma=32'd5;row=32'd298;
#400 gamma=32'd2;row=32'd198;
#400 gamma=32'd1;row=32'd256;
#400 gamma=32'd1;row=32'd397;
#400 gamma=32'd4;row=32'd212;
#400 gamma=32'd2;row=32'd500;
#400 gamma=32'd2;row=32'd440;
#400 gamma=32'd2;row=32'd101;
#400 gamma=32'd4;row=32'd520;
#400 gamma=32'd3;row=32'd93;
#400 gamma=32'd2;row=32'd388;
#400 gamma=32'd5;row=32'd52;
#400 gamma=32'd3;row=32'd103;
#400 gamma=32'd1;row=32'd298;
#400 gamma=32'd1;row=32'd185;
#400 gamma=32'd2;row=32'd248;
#400 gamma=32'd3;row=32'd329;
#400 gamma=32'd4;row=32'd137;
#400 gamma=32'd2;row=32'd289;
#400 gamma=32'd2;row=32'd358;
#400 gamma=32'd1;row=32'd67;
#400 gamma=32'd2;row=32'd42;
#400 gamma=32'd4;row=32'd217;
#400 gamma=32'd1;row=32'd290;
#400 gamma=32'd1;row=32'd119;
#400 gamma=32'd3;row=32'd406;
#400 gamma=32'd2;row=32'd343;
#400 gamma=32'd4;row=32'd147;
#400 gamma=32'd3;row=32'd559;
#400 gamma=32'd5;row=32'd295;
#400 gamma=32'd2;row=32'd332;
#400 gamma=32'd5;row=32'd247;
#400 gamma=32'd3;row=32'd304;
#400 gamma=32'd3;row=32'd267;
#400 gamma=32'd4;row=32'd509;
#400 gamma=32'd1;row=32'd4;
#400 gamma=32'd2;row=32'd187;
#400 gamma=32'd2;row=32'd365;
#400 gamma=32'd4;row=32'd551;
#400 gamma=32'd3;row=32'd197;
#400 gamma=32'd2;row=32'd416;
#400 gamma=32'd2;row=32'd63;
#400 gamma=32'd4;row=32'd253;
#400 gamma=32'd2;row=32'd120;
#400 gamma=32'd5;row=32'd393;
#400 gamma=32'd5;row=32'd535;
#400 gamma=32'd4;row=32'd199;
#400 gamma=32'd3;row=32'd181;
#400 gamma=32'd3;row=32'd419;
#400 gamma=32'd2;row=32'd65;
#400 gamma=32'd3;row=32'd487;
#400 gamma=32'd5;row=32'd432;
#400 gamma=32'd3;row=32'd215;
#400 gamma=32'd4;row=32'd211;
#400 gamma=32'd1;row=32'd265;
#400 gamma=32'd2;row=32'd8;
#400 gamma=32'd1;row=32'd376;
#400 gamma=32'd2;row=32'd0;
#400 gamma=32'd2;row=32'd535;
#400 gamma=32'd5;row=32'd109;
#400 gamma=32'd4;row=32'd233;
#400 gamma=32'd3;row=32'd530;
#400 gamma=32'd1;row=32'd477;
#400 gamma=32'd3;row=32'd302;
#400 gamma=32'd2;row=32'd381;
#400 gamma=32'd1;row=32'd203;
#400 gamma=32'd4;row=32'd138;
#400 gamma=32'd5;row=32'd143;
#400 gamma=32'd1;row=32'd98;
#400 gamma=32'd4;row=32'd71;
#400 gamma=32'd1;row=32'd126;
#400 gamma=32'd5;row=32'd245;
#400 gamma=32'd2;row=32'd109;
#400 gamma=32'd5;row=32'd6;
#400 gamma=32'd5;row=32'd223;
#400 gamma=32'd4;row=32'd155;
#400 gamma=32'd2;row=32'd145;
#400 gamma=32'd3;row=32'd501;
#400 gamma=32'd5;row=32'd294;
#400 gamma=32'd5;row=32'd494;
#400 gamma=32'd1;row=32'd289;
#400 gamma=32'd4;row=32'd341;
#400 gamma=32'd2;row=32'd257;
#400 gamma=32'd4;row=32'd442;
#400 gamma=32'd3;row=32'd12;
#400 gamma=32'd2;row=32'd71;
#400 gamma=32'd2;row=32'd505;
#400 gamma=32'd2;row=32'd332;
#400 gamma=32'd3;row=32'd138;
#400 gamma=32'd3;row=32'd304;
#400 gamma=32'd1;row=32'd541;
#400 gamma=32'd3;row=32'd241;
#400 gamma=32'd3;row=32'd228;
#400 gamma=32'd5;row=32'd86;
#400 gamma=32'd5;row=32'd232;
#400 gamma=32'd5;row=32'd392;
#400 gamma=32'd1;row=32'd282;
#400 gamma=32'd2;row=32'd477;
#400 gamma=32'd2;row=32'd328;
#400 gamma=32'd5;row=32'd312;
#400 gamma=32'd1;row=32'd215;
#400 gamma=32'd5;row=32'd111;
#400 gamma=32'd5;row=32'd324;
#400 gamma=32'd2;row=32'd477;
#400 gamma=32'd4;row=32'd531;
#400 gamma=32'd4;row=32'd482;
#400 gamma=32'd3;row=32'd283;
#400 gamma=32'd5;row=32'd423;
#400 gamma=32'd5;row=32'd366;
#400 gamma=32'd5;row=32'd28;
#400 gamma=32'd2;row=32'd407;
#400 gamma=32'd4;row=32'd230;
#400 gamma=32'd1;row=32'd135;
#400 gamma=32'd1;row=32'd183;
#400 gamma=32'd1;row=32'd131;
#400 gamma=32'd5;row=32'd173;
#400 gamma=32'd5;row=32'd161;
#400 gamma=32'd3;row=32'd116;
#400 gamma=32'd4;row=32'd544;
#400 gamma=32'd5;row=32'd121;
#400 gamma=32'd1;row=32'd546;
#400 gamma=32'd1;row=32'd258;
#400 gamma=32'd3;row=32'd510;
#400 gamma=32'd5;row=32'd21;
#400 gamma=32'd5;row=32'd362;
#400 gamma=32'd3;row=32'd99;
#400 gamma=32'd5;row=32'd146;
#400 gamma=32'd2;row=32'd94;
#400 gamma=32'd2;row=32'd399;
#400 gamma=32'd2;row=32'd218;
#400 gamma=32'd1;row=32'd315;
#400 gamma=32'd4;row=32'd244;
#400 gamma=32'd2;row=32'd72;
#400 gamma=32'd2;row=32'd391;
#400 gamma=32'd2;row=32'd213;
#400 gamma=32'd4;row=32'd312;
#400 gamma=32'd4;row=32'd235;
#400 gamma=32'd1;row=32'd154;
#400 gamma=32'd3;row=32'd149;
#400 gamma=32'd1;row=32'd414;
#400 gamma=32'd3;row=32'd287;
#400 gamma=32'd4;row=32'd53;
#400 gamma=32'd5;row=32'd339;
#400 gamma=32'd5;row=32'd372;
#400 gamma=32'd3;row=32'd455;
#400 gamma=32'd2;row=32'd277;
#400 gamma=32'd4;row=32'd37;
#400 gamma=32'd5;row=32'd14;
#400 gamma=32'd5;row=32'd326;
#400 gamma=32'd5;row=32'd263;
#400 gamma=32'd1;row=32'd508;
#400 gamma=32'd3;row=32'd505;
#400 gamma=32'd4;row=32'd212;
#400 gamma=32'd2;row=32'd429;
#400 gamma=32'd2;row=32'd292;
#400 gamma=32'd4;row=32'd515;
#400 gamma=32'd2;row=32'd313;
#400 gamma=32'd5;row=32'd440;
#400 gamma=32'd4;row=32'd389;
#400 gamma=32'd2;row=32'd215;
#400 gamma=32'd5;row=32'd33;
#400 gamma=32'd1;row=32'd344;
#400 gamma=32'd5;row=32'd135;
#400 gamma=32'd2;row=32'd113;
#400 gamma=32'd3;row=32'd314;
#400 gamma=32'd5;row=32'd22;
#400 gamma=32'd1;row=32'd326;
#400 gamma=32'd5;row=32'd498;
#400 gamma=32'd5;row=32'd545;
#400 gamma=32'd5;row=32'd32;
#400 gamma=32'd4;row=32'd347;
#400 gamma=32'd4;row=32'd381;
#400 gamma=32'd3;row=32'd435;
#400 gamma=32'd2;row=32'd420;
#400 gamma=32'd2;row=32'd101;
#400 gamma=32'd1;row=32'd303;
#400 gamma=32'd4;row=32'd64;
#400 gamma=32'd4;row=32'd244;
#400 gamma=32'd5;row=32'd429;
#400 gamma=32'd4;row=32'd406;
#400 gamma=32'd5;row=32'd172;
#400 gamma=32'd1;row=32'd500;
#400 gamma=32'd1;row=32'd36;
#400 gamma=32'd2;row=32'd282;
#400 gamma=32'd1;row=32'd456;
#400 gamma=32'd4;row=32'd426;
#400 gamma=32'd1;row=32'd126;
#400 gamma=32'd1;row=32'd68;
#400 gamma=32'd1;row=32'd362;
#400 gamma=32'd1;row=32'd394;
#400 gamma=32'd2;row=32'd541;
#400 gamma=32'd4;row=32'd322;
#400 gamma=32'd2;row=32'd541;
#400 gamma=32'd1;row=32'd88;
#400 gamma=32'd2;row=32'd175;
#400 gamma=32'd3;row=32'd501;
#400 gamma=32'd4;row=32'd79;
#400 gamma=32'd1;row=32'd52;
#400 gamma=32'd3;row=32'd396;
#400 gamma=32'd2;row=32'd174;
#400 gamma=32'd3;row=32'd14;
#400 gamma=32'd2;row=32'd40;
#400 gamma=32'd5;row=32'd435;
#400 gamma=32'd2;row=32'd28;
#400 gamma=32'd1;row=32'd443;
#400 gamma=32'd1;row=32'd466;
#400 gamma=32'd2;row=32'd155;
#400 gamma=32'd5;row=32'd472;
#400 gamma=32'd2;row=32'd75;
#400 gamma=32'd1;row=32'd506;
#400 gamma=32'd3;row=32'd217;
#400 gamma=32'd4;row=32'd448;
#400 gamma=32'd4;row=32'd296;
#400 gamma=32'd3;row=32'd142;
#400 gamma=32'd4;row=32'd160;
#400 gamma=32'd2;row=32'd95;
#400 gamma=32'd2;row=32'd111;
#400 gamma=32'd2;row=32'd46;
#400 gamma=32'd1;row=32'd342;
#400 gamma=32'd2;row=32'd461;
#400 gamma=32'd2;row=32'd43;
#400 gamma=32'd5;row=32'd265;
#400 gamma=32'd3;row=32'd481;
#400 gamma=32'd3;row=32'd159;
#400 gamma=32'd4;row=32'd101;
#400 gamma=32'd2;row=32'd473;
#400 gamma=32'd1;row=32'd479;
#400 gamma=32'd1;row=32'd461;
#400 gamma=32'd3;row=32'd465;
#400 gamma=32'd4;row=32'd425;
#400 gamma=32'd5;row=32'd508;
#400 gamma=32'd3;row=32'd311;
#400 gamma=32'd3;row=32'd89;
#400 gamma=32'd3;row=32'd328;
#400 gamma=32'd5;row=32'd281;
#400 gamma=32'd2;row=32'd316;
#400 gamma=32'd4;row=32'd116;
#400 gamma=32'd3;row=32'd342;
#400 gamma=32'd1;row=32'd332;
#400 gamma=32'd5;row=32'd162;
#400 gamma=32'd1;row=32'd219;
#400 gamma=32'd5;row=32'd205;
#400 gamma=32'd3;row=32'd57;
#400 gamma=32'd5;row=32'd13;
#400 gamma=32'd1;row=32'd111;
#400 gamma=32'd3;row=32'd112;
#400 gamma=32'd1;row=32'd233;
#400 gamma=32'd1;row=32'd137;
#400 gamma=32'd4;row=32'd147;
#400 gamma=32'd2;row=32'd465;
#400 gamma=32'd3;row=32'd113;
#400 gamma=32'd5;row=32'd549;
#400 gamma=32'd1;row=32'd104;
#400 gamma=32'd1;row=32'd477;
#400 gamma=32'd1;row=32'd468;
#400 gamma=32'd2;row=32'd388;
#400 gamma=32'd2;row=32'd395;
#400 gamma=32'd4;row=32'd253;
#400 gamma=32'd1;row=32'd267;
#400 gamma=32'd4;row=32'd433;
#400 gamma=32'd3;row=32'd477;
#400 gamma=32'd2;row=32'd436;
#400 gamma=32'd1;row=32'd322;
#400 gamma=32'd1;row=32'd421;
#400 gamma=32'd1;row=32'd98;
#400 gamma=32'd5;row=32'd197;
#400 gamma=32'd2;row=32'd489;
#400 gamma=32'd5;row=32'd101;
#400 gamma=32'd4;row=32'd453;
#400 gamma=32'd1;row=32'd260;
#400 gamma=32'd2;row=32'd4;
#400 gamma=32'd5;row=32'd464;
#400 gamma=32'd2;row=32'd252;
#400 gamma=32'd2;row=32'd231;
#400 gamma=32'd1;row=32'd48;
#400 gamma=32'd2;row=32'd544;
#400 gamma=32'd3;row=32'd340;
#400 gamma=32'd5;row=32'd176;
#400 gamma=32'd1;row=32'd449;
#400 gamma=32'd3;row=32'd30;
#400 gamma=32'd5;row=32'd477;
#400 gamma=32'd1;row=32'd150;
#400 gamma=32'd5;row=32'd530;
#400 gamma=32'd1;row=32'd456;
#400 gamma=32'd1;row=32'd231;
#400 gamma=32'd2;row=32'd158;
#400 gamma=32'd2;row=32'd386;
#400 gamma=32'd4;row=32'd298;
#400 gamma=32'd5;row=32'd79;
#400 gamma=32'd3;row=32'd515;
#400 gamma=32'd4;row=32'd484;
#400 gamma=32'd3;row=32'd219;
#400 gamma=32'd3;row=32'd83;
#400 gamma=32'd4;row=32'd174;
#400 gamma=32'd4;row=32'd130;
#400 gamma=32'd4;row=32'd411;
#400 gamma=32'd5;row=32'd435;
#400 gamma=32'd4;row=32'd227;
#400 gamma=32'd4;row=32'd219;
#400 gamma=32'd5;row=32'd235;
#400 gamma=32'd3;row=32'd556;
#400 gamma=32'd4;row=32'd131;
#400 gamma=32'd2;row=32'd70;
#400 gamma=32'd4;row=32'd116;
#400 gamma=32'd2;row=32'd49;
#400 gamma=32'd4;row=32'd106;
#400 gamma=32'd5;row=32'd129;
#400 gamma=32'd1;row=32'd91;
#400 gamma=32'd4;row=32'd176;
#400 gamma=32'd5;row=32'd273;
#400 gamma=32'd3;row=32'd305;
#400 gamma=32'd4;row=32'd469;
#400 gamma=32'd4;row=32'd233;
#400 gamma=32'd2;row=32'd477;
#400 gamma=32'd1;row=32'd528;
#400 gamma=32'd1;row=32'd58;
#400 gamma=32'd2;row=32'd87;
#400 gamma=32'd5;row=32'd464;
#400 gamma=32'd4;row=32'd81;
#400 gamma=32'd3;row=32'd429;
#400 gamma=32'd3;row=32'd467;
#400 gamma=32'd5;row=32'd497;
#400 gamma=32'd1;row=32'd345;
#400 gamma=32'd2;row=32'd433;
#400 gamma=32'd3;row=32'd296;
#400 gamma=32'd4;row=32'd22;
#400 gamma=32'd1;row=32'd503;
#400 gamma=32'd5;row=32'd306;
#400 gamma=32'd1;row=32'd341;
#400 gamma=32'd2;row=32'd36;
#400 gamma=32'd4;row=32'd524;
#400 gamma=32'd3;row=32'd221;
#400 gamma=32'd3;row=32'd485;
#400 gamma=32'd2;row=32'd472;
#400 gamma=32'd3;row=32'd417;
#400 gamma=32'd4;row=32'd353;
#400 gamma=32'd3;row=32'd295;
#400 gamma=32'd1;row=32'd276;
#400 gamma=32'd3;row=32'd526;
#400 gamma=32'd3;row=32'd6;
#400 gamma=32'd4;row=32'd215;
#400 gamma=32'd2;row=32'd267;
#400 gamma=32'd5;row=32'd364;
#400 gamma=32'd1;row=32'd279;
#400 gamma=32'd2;row=32'd276;
#400 gamma=32'd5;row=32'd98;
#400 gamma=32'd1;row=32'd540;
#400 gamma=32'd5;row=32'd253;
#400 gamma=32'd1;row=32'd198;
#400 gamma=32'd1;row=32'd304;
#400 gamma=32'd2;row=32'd364;
#400 gamma=32'd1;row=32'd286;
#400 gamma=32'd3;row=32'd29;
#400 gamma=32'd1;row=32'd99;
#400 gamma=32'd4;row=32'd156;
#400 gamma=32'd3;row=32'd337;
#400 gamma=32'd4;row=32'd83;
#400 gamma=32'd2;row=32'd528;
#400 gamma=32'd4;row=32'd110;
#400 gamma=32'd4;row=32'd224;
#400 gamma=32'd4;row=32'd292;
#400 gamma=32'd5;row=32'd451;
#400 gamma=32'd5;row=32'd251;
#400 gamma=32'd5;row=32'd1;
#400 gamma=32'd2;row=32'd278;
#400 gamma=32'd4;row=32'd108;
#400 gamma=32'd4;row=32'd552;
#400 gamma=32'd2;row=32'd503;
#400 gamma=32'd3;row=32'd496;
#400 gamma=32'd1;row=32'd60;
#400 gamma=32'd3;row=32'd224;
#400 gamma=32'd4;row=32'd438;
#400 gamma=32'd4;row=32'd428;
#400 gamma=32'd3;row=32'd34;
#400 gamma=32'd1;row=32'd232;
#400 gamma=32'd4;row=32'd108;
#400 gamma=32'd5;row=32'd2;
#400 gamma=32'd3;row=32'd51;
#400 gamma=32'd3;row=32'd436;
#400 gamma=32'd4;row=32'd442;
#400 gamma=32'd1;row=32'd428;
#400 gamma=32'd1;row=32'd153;
#400 gamma=32'd1;row=32'd161;
#400 gamma=32'd3;row=32'd394;
#400 gamma=32'd2;row=32'd212;
#400 gamma=32'd2;row=32'd499;
#400 gamma=32'd3;row=32'd274;
#400 gamma=32'd4;row=32'd368;
#400 gamma=32'd3;row=32'd299;
#400 gamma=32'd2;row=32'd359;
#400 gamma=32'd2;row=32'd105;
#400 gamma=32'd1;row=32'd369;
#400 gamma=32'd2;row=32'd84;
#400 gamma=32'd4;row=32'd147;
#400 gamma=32'd5;row=32'd221;
#400 gamma=32'd3;row=32'd477;
#400 gamma=32'd1;row=32'd523;
#400 gamma=32'd4;row=32'd555;
#400 gamma=32'd2;row=32'd519;
#400 gamma=32'd5;row=32'd208;
#400 gamma=32'd3;row=32'd468;
#400 gamma=32'd4;row=32'd407;
#400 gamma=32'd4;row=32'd350;
#400 gamma=32'd3;row=32'd234;
#400 gamma=32'd3;row=32'd360;
#400 gamma=32'd1;row=32'd277;
#400 gamma=32'd2;row=32'd357;
#400 gamma=32'd3;row=32'd159;
#400 gamma=32'd1;row=32'd278;
#400 gamma=32'd1;row=32'd175;
#400 gamma=32'd5;row=32'd361;
#400 gamma=32'd2;row=32'd195;
#400 gamma=32'd5;row=32'd344;
#400 gamma=32'd2;row=32'd548;
#400 gamma=32'd1;row=32'd231;
#400 gamma=32'd1;row=32'd546;
#400 gamma=32'd2;row=32'd297;
#400 gamma=32'd5;row=32'd37;
#400 gamma=32'd3;row=32'd349;
#400 gamma=32'd1;row=32'd141;
#400 gamma=32'd4;row=32'd435;
#400 gamma=32'd3;row=32'd28;
#400 gamma=32'd2;row=32'd67;
#400 gamma=32'd1;row=32'd184;
#400 gamma=32'd4;row=32'd200;
#400 gamma=32'd2;row=32'd238;
#400 gamma=32'd4;row=32'd216;
#400 gamma=32'd3;row=32'd234;
#400 gamma=32'd2;row=32'd487;
#400 gamma=32'd1;row=32'd531;
#400 gamma=32'd2;row=32'd146;
#400 gamma=32'd1;row=32'd396;
#400 gamma=32'd2;row=32'd541;
#400 gamma=32'd3;row=32'd322;
#400 gamma=32'd3;row=32'd92;
#400 gamma=32'd2;row=32'd492;
#400 gamma=32'd5;row=32'd24;
#400 gamma=32'd3;row=32'd272;
#400 gamma=32'd3;row=32'd0;
#400 gamma=32'd2;row=32'd455;
#400 gamma=32'd5;row=32'd56;
#400 gamma=32'd1;row=32'd532;
#400 gamma=32'd2;row=32'd213;
#400 gamma=32'd2;row=32'd69;
#400 gamma=32'd4;row=32'd321;
#400 gamma=32'd2;row=32'd527;
#400 gamma=32'd3;row=32'd547;
#400 gamma=32'd3;row=32'd89;
#400 gamma=32'd4;row=32'd548;
#400 gamma=32'd5;row=32'd34;
#400 gamma=32'd1;row=32'd316;
#400 gamma=32'd1;row=32'd291;
#400 gamma=32'd2;row=32'd121;
#400 gamma=32'd5;row=32'd84;
#400 gamma=32'd1;row=32'd102;
#400 gamma=32'd5;row=32'd203;
#400 gamma=32'd1;row=32'd148;
#400 gamma=32'd2;row=32'd142;
#400 gamma=32'd5;row=32'd94;
#400 gamma=32'd3;row=32'd241;
#400 gamma=32'd2;row=32'd367;
#400 gamma=32'd4;row=32'd331;
#400 gamma=32'd1;row=32'd213;
#400 gamma=32'd5;row=32'd94;
#400 gamma=32'd5;row=32'd404;
#400 gamma=32'd2;row=32'd199;
#400 gamma=32'd3;row=32'd162;
#400 gamma=32'd1;row=32'd323;
#400 gamma=32'd2;row=32'd264;
#400 gamma=32'd5;row=32'd114;
#400 gamma=32'd1;row=32'd390;
#400 gamma=32'd3;row=32'd346;
#400 gamma=32'd5;row=32'd469;
#400 gamma=32'd2;row=32'd79;
#400 gamma=32'd3;row=32'd31;
#400 gamma=32'd4;row=32'd411;
#400 gamma=32'd5;row=32'd554;
#400 gamma=32'd5;row=32'd474;
#400 gamma=32'd3;row=32'd387;
#400 gamma=32'd3;row=32'd452;
#400 gamma=32'd3;row=32'd19;
#400 gamma=32'd4;row=32'd408;
#400 gamma=32'd4;row=32'd325;
#400 gamma=32'd4;row=32'd230;
#400 gamma=32'd5;row=32'd129;
#400 gamma=32'd1;row=32'd394;
#400 gamma=32'd5;row=32'd313;
#400 gamma=32'd2;row=32'd374;
#400 gamma=32'd3;row=32'd294;
#400 gamma=32'd2;row=32'd332;
#400 gamma=32'd3;row=32'd223;
#400 gamma=32'd4;row=32'd80;
#400 gamma=32'd4;row=32'd419;
#400 gamma=32'd4;row=32'd123;
#400 gamma=32'd3;row=32'd491;
#400 gamma=32'd3;row=32'd235;
#400 gamma=32'd5;row=32'd440;
#400 gamma=32'd3;row=32'd345;
#400 gamma=32'd5;row=32'd47;
#400 gamma=32'd3;row=32'd237;
#400 gamma=32'd3;row=32'd176;
#400 gamma=32'd4;row=32'd415;
#400 gamma=32'd1;row=32'd423;
#400 gamma=32'd2;row=32'd215;
#400 gamma=32'd2;row=32'd17;
#400 gamma=32'd1;row=32'd296;
#400 gamma=32'd4;row=32'd104;
#400 gamma=32'd2;row=32'd521;
#400 gamma=32'd2;row=32'd62;
#400 gamma=32'd2;row=32'd307;
#400 gamma=32'd1;row=32'd479;
#400 gamma=32'd3;row=32'd330;
#400 gamma=32'd3;row=32'd313;
#400 gamma=32'd3;row=32'd14;
#400 gamma=32'd1;row=32'd93;
#400 gamma=32'd4;row=32'd193;
#400 gamma=32'd5;row=32'd157;
#400 gamma=32'd2;row=32'd480;
#400 gamma=32'd5;row=32'd219;
#400 gamma=32'd4;row=32'd294;
#400 gamma=32'd3;row=32'd425;
#400 gamma=32'd2;row=32'd190;
#400 gamma=32'd5;row=32'd58;
#400 gamma=32'd1;row=32'd530;
#400 gamma=32'd3;row=32'd286;
#400 gamma=32'd5;row=32'd253;
#400 gamma=32'd2;row=32'd396;
#400 gamma=32'd4;row=32'd384;
#400 gamma=32'd2;row=32'd218;
#400 gamma=32'd3;row=32'd478;
#400 gamma=32'd5;row=32'd485;
#400 gamma=32'd4;row=32'd42;
#400 gamma=32'd1;row=32'd297;
#400 gamma=32'd3;row=32'd429;
#400 gamma=32'd5;row=32'd44;
#400 gamma=32'd1;row=32'd348;
#400 gamma=32'd1;row=32'd11;
#400 gamma=32'd2;row=32'd325;
#400 gamma=32'd1;row=32'd25;
#400 gamma=32'd1;row=32'd254;
#400 gamma=32'd3;row=32'd401;
#400 gamma=32'd5;row=32'd390;
#400 gamma=32'd3;row=32'd52;
#400 gamma=32'd2;row=32'd471;
#400 gamma=32'd1;row=32'd289;
#400 gamma=32'd4;row=32'd320;
#400 gamma=32'd5;row=32'd286;
#400 gamma=32'd4;row=32'd417;
#400 gamma=32'd1;row=32'd114;
#400 gamma=32'd3;row=32'd416;
#400 gamma=32'd4;row=32'd208;
#400 gamma=32'd5;row=32'd3;
#400 gamma=32'd2;row=32'd217;
#400 gamma=32'd1;row=32'd250;
#400 gamma=32'd2;row=32'd405;
#400 gamma=32'd4;row=32'd402;
#400 gamma=32'd4;row=32'd469;
#400 gamma=32'd2;row=32'd161;
#400 gamma=32'd4;row=32'd292;
#400 gamma=32'd5;row=32'd508;
#400 gamma=32'd5;row=32'd125;
#400 gamma=32'd2;row=32'd285;
#400 gamma=32'd2;row=32'd119;
#400 gamma=32'd5;row=32'd277;
#400 gamma=32'd3;row=32'd22;
#400 gamma=32'd2;row=32'd343;
#400 gamma=32'd2;row=32'd459;
#400 gamma=32'd2;row=32'd258;
#400 gamma=32'd2;row=32'd9;
#400 gamma=32'd4;row=32'd163;
#400 gamma=32'd3;row=32'd521;
#400 gamma=32'd3;row=32'd436;
#400 gamma=32'd1;row=32'd364;
#400 gamma=32'd5;row=32'd157;
#400 gamma=32'd2;row=32'd78;
#400 gamma=32'd5;row=32'd278;
#400 gamma=32'd1;row=32'd348;
#400 gamma=32'd3;row=32'd443;
#400 gamma=32'd2;row=32'd22;
#400 gamma=32'd2;row=32'd335;
#400 gamma=32'd4;row=32'd229;
#400 gamma=32'd1;row=32'd541;
#400 gamma=32'd2;row=32'd234;
#400 gamma=32'd4;row=32'd64;
#400 gamma=32'd4;row=32'd11;
#400 gamma=32'd1;row=32'd555;
#400 gamma=32'd2;row=32'd378;
#400 gamma=32'd3;row=32'd78;
#400 gamma=32'd3;row=32'd551;
#400 gamma=32'd5;row=32'd277;
#400 gamma=32'd1;row=32'd441;
#400 gamma=32'd2;row=32'd430;
#400 gamma=32'd5;row=32'd225;
#400 gamma=32'd2;row=32'd276;
#400 gamma=32'd5;row=32'd500;
#400 gamma=32'd2;row=32'd394;
#400 gamma=32'd4;row=32'd411;
#400 gamma=32'd3;row=32'd464;
#400 gamma=32'd2;row=32'd56;
#400 gamma=32'd3;row=32'd544;
#400 gamma=32'd2;row=32'd491;
#400 gamma=32'd5;row=32'd74;
#400 gamma=32'd3;row=32'd296;
#400 gamma=32'd3;row=32'd86;
#400 gamma=32'd5;row=32'd138;
#400 gamma=32'd2;row=32'd380;
#400 gamma=32'd2;row=32'd35;
#400 gamma=32'd3;row=32'd211;
#400 gamma=32'd2;row=32'd365;
#400 gamma=32'd5;row=32'd291;
#400 gamma=32'd2;row=32'd33;
#400 gamma=32'd3;row=32'd418;
#400 gamma=32'd1;row=32'd223;
#400 gamma=32'd3;row=32'd485;
#400 gamma=32'd5;row=32'd530;
#400 gamma=32'd4;row=32'd436;
#400 gamma=32'd5;row=32'd323;
#400 gamma=32'd4;row=32'd460;
#400 gamma=32'd4;row=32'd63;
#400 gamma=32'd1;row=32'd257;
#400 gamma=32'd5;row=32'd95;
#400 gamma=32'd3;row=32'd294;
#400 gamma=32'd5;row=32'd13;
#400 gamma=32'd4;row=32'd429;
#400 gamma=32'd2;row=32'd38;
#400 gamma=32'd2;row=32'd48;
#400 gamma=32'd2;row=32'd72;
#400 gamma=32'd1;row=32'd209;
#400 gamma=32'd1;row=32'd15;
#400 gamma=32'd2;row=32'd426;
#400 gamma=32'd2;row=32'd164;
#400 gamma=32'd3;row=32'd157;
#400 gamma=32'd5;row=32'd546;
#400 gamma=32'd2;row=32'd393;
#400 gamma=32'd3;row=32'd159;
#400 gamma=32'd3;row=32'd93;
#400 gamma=32'd5;row=32'd74;
#400 gamma=32'd2;row=32'd40;
#400 gamma=32'd5;row=32'd327;
#400 gamma=32'd1;row=32'd447;
#400 gamma=32'd2;row=32'd482;
#400 gamma=32'd5;row=32'd559;
#400 gamma=32'd4;row=32'd8;
#400 gamma=32'd4;row=32'd284;
#400 gamma=32'd2;row=32'd220;
#400 gamma=32'd2;row=32'd65;
#400 gamma=32'd3;row=32'd344;
#400 gamma=32'd5;row=32'd117;
#400 gamma=32'd2;row=32'd110;
#400 gamma=32'd5;row=32'd253;
#400 gamma=32'd4;row=32'd548;
#400 gamma=32'd3;row=32'd454;
#400 gamma=32'd5;row=32'd170;
#400 gamma=32'd3;row=32'd99;
#400 gamma=32'd5;row=32'd10;
#400 gamma=32'd5;row=32'd120;
#400 gamma=32'd4;row=32'd355;
#400 gamma=32'd5;row=32'd244;
#400 gamma=32'd5;row=32'd17;
#400 gamma=32'd4;row=32'd9;
#400 gamma=32'd1;row=32'd2;
#400 gamma=32'd3;row=32'd142;
#400 gamma=32'd3;row=32'd35;
#400 gamma=32'd5;row=32'd204;
#400 gamma=32'd2;row=32'd132;
#400 gamma=32'd2;row=32'd93;
#400 gamma=32'd5;row=32'd115;
#400 gamma=32'd5;row=32'd202;
#400 gamma=32'd5;row=32'd301;
#400 gamma=32'd2;row=32'd182;
#400 gamma=32'd2;row=32'd76;
#400 gamma=32'd5;row=32'd458;
#400 gamma=32'd1;row=32'd552;
#400 gamma=32'd1;row=32'd330;
#400 gamma=32'd2;row=32'd201;
#400 gamma=32'd3;row=32'd222;
#400 gamma=32'd3;row=32'd417;
#400 gamma=32'd3;row=32'd319;
#400 gamma=32'd2;row=32'd151;
#400 gamma=32'd5;row=32'd354;
#400 gamma=32'd1;row=32'd544;
#400 gamma=32'd2;row=32'd81;
#400 gamma=32'd5;row=32'd175;
#400 gamma=32'd2;row=32'd70;
#400 gamma=32'd5;row=32'd243;
#400 gamma=32'd5;row=32'd205;
#400 gamma=32'd1;row=32'd23;
#400 gamma=32'd1;row=32'd547;
#400 gamma=32'd4;row=32'd416;
#400 gamma=32'd5;row=32'd405;
#400 gamma=32'd5;row=32'd524;
#400 gamma=32'd5;row=32'd351;
#400 gamma=32'd5;row=32'd433;
#400 gamma=32'd3;row=32'd376;
#400 gamma=32'd3;row=32'd129;
#400 gamma=32'd1;row=32'd32;
#400 gamma=32'd3;row=32'd478;
#400 gamma=32'd2;row=32'd451;
#400 gamma=32'd5;row=32'd377;
#400 gamma=32'd1;row=32'd330;
#400 gamma=32'd1;row=32'd242;
#400 gamma=32'd3;row=32'd544;
#400 gamma=32'd1;row=32'd390;
#400 gamma=32'd3;row=32'd144;
#400 gamma=32'd1;row=32'd274;
#400 gamma=32'd5;row=32'd143;
#400 gamma=32'd4;row=32'd97;
#400 gamma=32'd3;row=32'd471;
#400 gamma=32'd1;row=32'd172;
#400 gamma=32'd5;row=32'd426;
#400 gamma=32'd4;row=32'd2;
#400 gamma=32'd1;row=32'd507;
#400 gamma=32'd5;row=32'd494;
#400 gamma=32'd3;row=32'd272;
#400 gamma=32'd1;row=32'd39;
#400 gamma=32'd3;row=32'd507;
#400 gamma=32'd5;row=32'd394;
#400 gamma=32'd5;row=32'd136;
#400 gamma=32'd5;row=32'd72;
#400 gamma=32'd1;row=32'd524;
#400 gamma=32'd3;row=32'd249;
#400 gamma=32'd1;row=32'd531;
#400 gamma=32'd1;row=32'd330;
#400 gamma=32'd2;row=32'd219;
#400 gamma=32'd4;row=32'd456;
#400 gamma=32'd5;row=32'd511;
#400 gamma=32'd5;row=32'd399;
#400 gamma=32'd3;row=32'd312;
#400 gamma=32'd1;row=32'd338;
#400 gamma=32'd5;row=32'd375;
#400 gamma=32'd1;row=32'd18;
#400 gamma=32'd1;row=32'd78;
#400 gamma=32'd5;row=32'd104;
#400 gamma=32'd1;row=32'd209;
#400 gamma=32'd2;row=32'd519;
#400 gamma=32'd5;row=32'd98;
#400 gamma=32'd4;row=32'd544;
#400 gamma=32'd4;row=32'd16;
#400 gamma=32'd4;row=32'd462;
#400 gamma=32'd2;row=32'd321;
#400 gamma=32'd4;row=32'd397;
#400 gamma=32'd5;row=32'd192;
#400 gamma=32'd2;row=32'd415;
#400 gamma=32'd5;row=32'd526;
#400 gamma=32'd4;row=32'd528;
#400 gamma=32'd1;row=32'd120;
#400 gamma=32'd1;row=32'd557;
#400 gamma=32'd2;row=32'd309;
#400 gamma=32'd5;row=32'd26;
#400 gamma=32'd3;row=32'd319;
#400 gamma=32'd1;row=32'd74;
#400 gamma=32'd1;row=32'd83;
#400 gamma=32'd3;row=32'd264;
#400 gamma=32'd5;row=32'd460;
#400 gamma=32'd2;row=32'd224;
#400 gamma=32'd3;row=32'd31;
#400 gamma=32'd3;row=32'd252;
#400 gamma=32'd5;row=32'd392;
#400 gamma=32'd4;row=32'd499;
#400 gamma=32'd3;row=32'd445;
#400 gamma=32'd5;row=32'd8;
#400 gamma=32'd1;row=32'd215;
#400 gamma=32'd5;row=32'd503;
#400 gamma=32'd4;row=32'd389;
#400 gamma=32'd5;row=32'd484;
#400 gamma=32'd5;row=32'd445;
#400 gamma=32'd3;row=32'd25;
#400 gamma=32'd4;row=32'd30;
#400 gamma=32'd1;row=32'd172;
#400 gamma=32'd3;row=32'd280;
#400 gamma=32'd2;row=32'd95;
#400 gamma=32'd5;row=32'd210;
#400 gamma=32'd3;row=32'd276;
#400 gamma=32'd3;row=32'd493;
#400 gamma=32'd4;row=32'd353;
#400 gamma=32'd1;row=32'd534;
#400 gamma=32'd5;row=32'd467;
#400 gamma=32'd5;row=32'd121;
#400 gamma=32'd1;row=32'd459;
#400 gamma=32'd5;row=32'd400;
#400 gamma=32'd5;row=32'd12;
#400 gamma=32'd1;row=32'd508;
#400 gamma=32'd1;row=32'd375;
#400 gamma=32'd2;row=32'd82;
#400 gamma=32'd5;row=32'd273;
#400 gamma=32'd3;row=32'd248;
#400 gamma=32'd1;row=32'd142;
#400 gamma=32'd3;row=32'd14;
#400 gamma=32'd4;row=32'd324;
#400 gamma=32'd3;row=32'd329;
#400 gamma=32'd5;row=32'd399;
#400 gamma=32'd5;row=32'd444;
#400 gamma=32'd3;row=32'd488;
#400 gamma=32'd2;row=32'd146;
#400 gamma=32'd2;row=32'd69;
#400 gamma=32'd5;row=32'd11;
#400 gamma=32'd4;row=32'd356;
#400 gamma=32'd3;row=32'd122;
#400 gamma=32'd1;row=32'd353;
#400 gamma=32'd5;row=32'd273;
#400 gamma=32'd2;row=32'd47;
#400 gamma=32'd1;row=32'd137;
#400 gamma=32'd2;row=32'd149;
#400 gamma=32'd4;row=32'd220;
#400 gamma=32'd3;row=32'd109;
#400 gamma=32'd3;row=32'd277;
#400 gamma=32'd2;row=32'd255;
#400 gamma=32'd1;row=32'd120;
#400 gamma=32'd3;row=32'd190;
#400 gamma=32'd2;row=32'd525;
#400 gamma=32'd2;row=32'd421;
#400 gamma=32'd3;row=32'd122;
#400 gamma=32'd5;row=32'd344;
#400 gamma=32'd5;row=32'd409;
#400 gamma=32'd3;row=32'd17;
#400 gamma=32'd4;row=32'd96;
#400 gamma=32'd5;row=32'd312;
#400 gamma=32'd3;row=32'd323;
#400 gamma=32'd2;row=32'd52;
#400 gamma=32'd5;row=32'd416;
#400 gamma=32'd5;row=32'd453;
#400 gamma=32'd2;row=32'd63;
#400 gamma=32'd1;row=32'd4;
#400 gamma=32'd3;row=32'd87;
#400 gamma=32'd5;row=32'd98;
#400 gamma=32'd3;row=32'd356;
#400 gamma=32'd4;row=32'd382;
#400 gamma=32'd2;row=32'd433;
#400 gamma=32'd3;row=32'd524;
#400 gamma=32'd5;row=32'd185;
#400 gamma=32'd2;row=32'd5;
#400 gamma=32'd4;row=32'd429;
#400 gamma=32'd1;row=32'd273;
#400 gamma=32'd5;row=32'd484;
#400 gamma=32'd5;row=32'd140;
#400 gamma=32'd2;row=32'd187;
#400 gamma=32'd4;row=32'd172;
#400 gamma=32'd2;row=32'd545;
#400 gamma=32'd4;row=32'd140;
#400 gamma=32'd3;row=32'd510;
#400 gamma=32'd5;row=32'd127;
#400 gamma=32'd3;row=32'd474;
#400 gamma=32'd3;row=32'd143;
#400 gamma=32'd3;row=32'd317;
#400 gamma=32'd3;row=32'd15;
#400 gamma=32'd1;row=32'd93;
#400 gamma=32'd4;row=32'd418;
#400 gamma=32'd3;row=32'd486;
#400 gamma=32'd4;row=32'd248;
#400 gamma=32'd1;row=32'd263;
#400 gamma=32'd3;row=32'd144;
#400 gamma=32'd4;row=32'd10;
#400 gamma=32'd4;row=32'd443;
#400 gamma=32'd2;row=32'd170;
#400 gamma=32'd4;row=32'd85;
#400 gamma=32'd2;row=32'd395;
#400 gamma=32'd5;row=32'd406;
#400 gamma=32'd1;row=32'd200;
#400 gamma=32'd5;row=32'd559;
#400 gamma=32'd3;row=32'd103;
#400 gamma=32'd3;row=32'd254;
#400 gamma=32'd1;row=32'd422;
#400 gamma=32'd2;row=32'd54;
#400 gamma=32'd1;row=32'd356;
#400 gamma=32'd3;row=32'd264;
#400 gamma=32'd4;row=32'd124;
#400 gamma=32'd4;row=32'd347;
#400 gamma=32'd5;row=32'd236;
#400 gamma=32'd5;row=32'd404;
#400 gamma=32'd3;row=32'd375;
#400 gamma=32'd4;row=32'd329;
#400 gamma=32'd1;row=32'd177;
#400 gamma=32'd5;row=32'd396;
#400 gamma=32'd4;row=32'd140;
#400 gamma=32'd3;row=32'd238;
#400 gamma=32'd2;row=32'd49;
#400 gamma=32'd2;row=32'd208;
#400 gamma=32'd3;row=32'd511;
#400 gamma=32'd1;row=32'd541;
#400 gamma=32'd5;row=32'd371;
#400 gamma=32'd4;row=32'd267;
#400 gamma=32'd4;row=32'd458;
#400 gamma=32'd1;row=32'd555;
#400 gamma=32'd2;row=32'd496;
#400 gamma=32'd4;row=32'd118;
#400 gamma=32'd1;row=32'd466;
#400 gamma=32'd1;row=32'd275;
#400 gamma=32'd5;row=32'd51;
#400 gamma=32'd4;row=32'd437;
#400 gamma=32'd2;row=32'd76;
#400 gamma=32'd2;row=32'd368;
#400 gamma=32'd5;row=32'd517;
#400 gamma=32'd5;row=32'd91;
#400 gamma=32'd5;row=32'd377;
#400 gamma=32'd3;row=32'd133;
#400 gamma=32'd3;row=32'd268;
#400 gamma=32'd5;row=32'd31;
#400 gamma=32'd5;row=32'd263;
#400 gamma=32'd1;row=32'd287;
#400 gamma=32'd3;row=32'd236;
#400 gamma=32'd3;row=32'd130;
#400 gamma=32'd3;row=32'd303;
#400 gamma=32'd5;row=32'd428;
#400 gamma=32'd5;row=32'd540;
#400 gamma=32'd3;row=32'd165;
#400 gamma=32'd5;row=32'd544;
#400 gamma=32'd4;row=32'd411;
#400 gamma=32'd2;row=32'd96;
#400 gamma=32'd1;row=32'd160;
#400 gamma=32'd5;row=32'd475;
#400 gamma=32'd4;row=32'd288;
#400 gamma=32'd3;row=32'd71;
#400 gamma=32'd2;row=32'd134;
#400 gamma=32'd3;row=32'd389;
#400 gamma=32'd4;row=32'd362;
#400 gamma=32'd1;row=32'd358;
#400 gamma=32'd3;row=32'd111;
#400 gamma=32'd1;row=32'd138;
#400 gamma=32'd3;row=32'd105;
#400 gamma=32'd2;row=32'd164;
#400 gamma=32'd1;row=32'd381;
#400 gamma=32'd1;row=32'd69;
#400 gamma=32'd1;row=32'd52;
#400 gamma=32'd5;row=32'd348;
#400 gamma=32'd5;row=32'd344;
#400 gamma=32'd2;row=32'd271;
#400 gamma=32'd4;row=32'd541;
#400 gamma=32'd2;row=32'd406;
#400 gamma=32'd3;row=32'd345;
#400 gamma=32'd4;row=32'd239;
#400 gamma=32'd1;row=32'd171;
#400 gamma=32'd4;row=32'd26;
#400 gamma=32'd3;row=32'd336;
#400 gamma=32'd4;row=32'd111;
#400 gamma=32'd3;row=32'd315;
#400 gamma=32'd1;row=32'd245;
#400 gamma=32'd2;row=32'd539;
#400 gamma=32'd3;row=32'd176;
#400 gamma=32'd3;row=32'd20;
#400 gamma=32'd1;row=32'd181;
#400 gamma=32'd2;row=32'd195;
#400 gamma=32'd1;row=32'd77;
#400 gamma=32'd3;row=32'd307;
#400 gamma=32'd5;row=32'd203;
#400 gamma=32'd5;row=32'd128;
#400 gamma=32'd3;row=32'd359;
#400 gamma=32'd2;row=32'd136;
#400 gamma=32'd1;row=32'd255;
#400 gamma=32'd1;row=32'd329;
#400 gamma=32'd3;row=32'd117;
#400 gamma=32'd5;row=32'd527;
#400 gamma=32'd5;row=32'd67;
#400 gamma=32'd5;row=32'd207;
#400 gamma=32'd2;row=32'd378;
#400 gamma=32'd1;row=32'd291;
#400 gamma=32'd1;row=32'd197;
#400 gamma=32'd2;row=32'd63;
#400 gamma=32'd4;row=32'd123;
#400 gamma=32'd1;row=32'd413;
#400 gamma=32'd1;row=32'd440;
#400 gamma=32'd5;row=32'd144;
#400 gamma=32'd1;row=32'd403;
#400 gamma=32'd2;row=32'd44;
#400 gamma=32'd4;row=32'd461;
#400 gamma=32'd1;row=32'd502;
#400 gamma=32'd1;row=32'd100;
#400 gamma=32'd3;row=32'd308;
#400 gamma=32'd3;row=32'd383;
#400 gamma=32'd5;row=32'd504;
#400 gamma=32'd2;row=32'd298;
#400 gamma=32'd3;row=32'd258;
#400 gamma=32'd1;row=32'd327;
#400 gamma=32'd3;row=32'd514;
#400 gamma=32'd4;row=32'd46;
#400 gamma=32'd2;row=32'd159;
#400 gamma=32'd2;row=32'd402;
#400 gamma=32'd2;row=32'd493;
#400 gamma=32'd1;row=32'd297;
#400 gamma=32'd3;row=32'd424;
#400 gamma=32'd4;row=32'd545;
#400 gamma=32'd3;row=32'd558;
#400 gamma=32'd1;row=32'd395;
#400 gamma=32'd3;row=32'd526;
#400 gamma=32'd5;row=32'd377;
#400 gamma=32'd1;row=32'd466;
#400 gamma=32'd4;row=32'd308;
#400 gamma=32'd1;row=32'd218;
#400 gamma=32'd4;row=32'd413;
#400 gamma=32'd1;row=32'd109;
#400 gamma=32'd2;row=32'd187;
#400 gamma=32'd4;row=32'd395;
#400 gamma=32'd2;row=32'd189;
#400 gamma=32'd1;row=32'd391;
#400 gamma=32'd5;row=32'd438;
#400 gamma=32'd5;row=32'd389;
#400 gamma=32'd4;row=32'd356;
#400 gamma=32'd5;row=32'd507;
#400 gamma=32'd4;row=32'd257;
#400 gamma=32'd1;row=32'd539;
#400 gamma=32'd3;row=32'd388;
#400 gamma=32'd1;row=32'd434;
#400 gamma=32'd3;row=32'd74;
#400 gamma=32'd4;row=32'd44;
#400 gamma=32'd5;row=32'd159;
#400 gamma=32'd5;row=32'd248;
#400 gamma=32'd4;row=32'd330;
#400 gamma=32'd2;row=32'd187;
#400 gamma=32'd5;row=32'd113;
#400 gamma=32'd4;row=32'd150;
#400 gamma=32'd1;row=32'd428;
#400 gamma=32'd3;row=32'd468;
#400 gamma=32'd4;row=32'd292;
#400 gamma=32'd5;row=32'd103;
#400 gamma=32'd2;row=32'd419;
#400 gamma=32'd2;row=32'd467;
#400 gamma=32'd2;row=32'd385;
#400 gamma=32'd3;row=32'd364;
#400 gamma=32'd2;row=32'd518;
#400 gamma=32'd4;row=32'd355;
#400 gamma=32'd3;row=32'd395;
#400 gamma=32'd1;row=32'd480;
#400 gamma=32'd5;row=32'd264;
#400 gamma=32'd5;row=32'd26;
#400 gamma=32'd1;row=32'd534;
#400 gamma=32'd5;row=32'd239;
#400 gamma=32'd4;row=32'd133;
#400 gamma=32'd1;row=32'd364;
#400 gamma=32'd3;row=32'd270;
#400 gamma=32'd3;row=32'd175;
#400 gamma=32'd2;row=32'd149;
#400 gamma=32'd3;row=32'd539;
#400 gamma=32'd4;row=32'd363;
#400 gamma=32'd5;row=32'd66;
#400 gamma=32'd1;row=32'd262;
#400 gamma=32'd1;row=32'd526;
#400 gamma=32'd2;row=32'd367;
#400 gamma=32'd4;row=32'd379;
#400 gamma=32'd5;row=32'd197;
#400 gamma=32'd4;row=32'd108;
#400 gamma=32'd4;row=32'd13;
#400 gamma=32'd1;row=32'd538;
#400 gamma=32'd4;row=32'd266;
#400 gamma=32'd5;row=32'd98;
#400 gamma=32'd3;row=32'd120;
#400 gamma=32'd1;row=32'd96;
#400 gamma=32'd1;row=32'd489;
#400 gamma=32'd1;row=32'd40;
#400 gamma=32'd2;row=32'd321;
#400 gamma=32'd2;row=32'd344;
#400 gamma=32'd4;row=32'd412;
#400 gamma=32'd3;row=32'd63;
#400 gamma=32'd4;row=32'd45;
#400 gamma=32'd3;row=32'd243;
#400 gamma=32'd5;row=32'd327;
#400 gamma=32'd5;row=32'd442;
#400 gamma=32'd2;row=32'd341;
#400 gamma=32'd3;row=32'd365;
#400 gamma=32'd5;row=32'd80;
#400 gamma=32'd5;row=32'd433;
#400 gamma=32'd1;row=32'd554;
#400 gamma=32'd1;row=32'd272;
#400 gamma=32'd5;row=32'd447;
#400 gamma=32'd1;row=32'd475;
#400 gamma=32'd3;row=32'd502;
#400 gamma=32'd5;row=32'd163;
#400 gamma=32'd3;row=32'd558;
#400 gamma=32'd4;row=32'd231;
#400 gamma=32'd1;row=32'd256;
#400 gamma=32'd5;row=32'd288;
#400 gamma=32'd4;row=32'd276;
#400 gamma=32'd2;row=32'd532;
#400 gamma=32'd4;row=32'd470;
#400 gamma=32'd3;row=32'd540;
#400 gamma=32'd1;row=32'd211;
#400 gamma=32'd3;row=32'd78;
#400 gamma=32'd5;row=32'd172;
#400 gamma=32'd5;row=32'd7;
#400 gamma=32'd3;row=32'd6;
#400 gamma=32'd2;row=32'd291;
#400 gamma=32'd4;row=32'd331;
#400 gamma=32'd5;row=32'd478;
#400 gamma=32'd4;row=32'd52;
#400 gamma=32'd2;row=32'd513;
#400 gamma=32'd1;row=32'd361;
#400 gamma=32'd5;row=32'd291;
#400 gamma=32'd1;row=32'd510;
#400 gamma=32'd1;row=32'd491;
#400 gamma=32'd2;row=32'd546;
#400 gamma=32'd2;row=32'd91;
#400 gamma=32'd1;row=32'd243;
#400 gamma=32'd1;row=32'd437;
#400 gamma=32'd5;row=32'd132;
#400 gamma=32'd4;row=32'd208;
#400 gamma=32'd2;row=32'd267;
#400 gamma=32'd3;row=32'd69;
#400 gamma=32'd5;row=32'd557;
#400 gamma=32'd1;row=32'd240;
#400 gamma=32'd3;row=32'd350;
#400 gamma=32'd2;row=32'd526;
#400 gamma=32'd5;row=32'd286;
#400 gamma=32'd4;row=32'd236;
#400 gamma=32'd4;row=32'd524;
#400 gamma=32'd3;row=32'd152;
#400 gamma=32'd5;row=32'd472;
#400 gamma=32'd5;row=32'd34;
#400 gamma=32'd1;row=32'd381;
#400 gamma=32'd3;row=32'd509;
#400 gamma=32'd3;row=32'd60;
#400 gamma=32'd2;row=32'd15;
#400 gamma=32'd1;row=32'd166;
#400 gamma=32'd4;row=32'd511;
#400 gamma=32'd4;row=32'd393;
#400 gamma=32'd3;row=32'd75;
#400 gamma=32'd1;row=32'd400;
#400 gamma=32'd2;row=32'd75;
#400 gamma=32'd5;row=32'd483;
#400 gamma=32'd5;row=32'd242;
#400 gamma=32'd2;row=32'd224;
#400 gamma=32'd1;row=32'd278;
#400 gamma=32'd1;row=32'd4;
#400 gamma=32'd2;row=32'd23;
#400 gamma=32'd3;row=32'd29;
#400 gamma=32'd1;row=32'd16;
#400 gamma=32'd4;row=32'd545;
#400 gamma=32'd3;row=32'd535;
#400 gamma=32'd1;row=32'd99;
#400 gamma=32'd2;row=32'd270;
#400 gamma=32'd1;row=32'd348;
#400 gamma=32'd1;row=32'd362;
#400 gamma=32'd4;row=32'd296;
#400 gamma=32'd3;row=32'd16;
#400 gamma=32'd2;row=32'd276;
#400 gamma=32'd3;row=32'd64;
#400 gamma=32'd3;row=32'd42;
#400 gamma=32'd3;row=32'd177;
#400 gamma=32'd1;row=32'd136;
#400 gamma=32'd1;row=32'd379;
#400 gamma=32'd1;row=32'd299;
#400 gamma=32'd2;row=32'd393;
#400 gamma=32'd1;row=32'd549;
#400 gamma=32'd4;row=32'd94;
#400 gamma=32'd3;row=32'd476;
#400 gamma=32'd1;row=32'd117;
#400 gamma=32'd2;row=32'd459;
#400 gamma=32'd5;row=32'd23;
#400 gamma=32'd1;row=32'd499;
#400 gamma=32'd4;row=32'd105;
#400 gamma=32'd2;row=32'd355;
#400 gamma=32'd5;row=32'd396;
#400 gamma=32'd1;row=32'd100;
#400 gamma=32'd1;row=32'd203;
#400 gamma=32'd4;row=32'd530;
#400 gamma=32'd5;row=32'd322;
#400 gamma=32'd4;row=32'd345;
#400 gamma=32'd5;row=32'd453;
#400 gamma=32'd3;row=32'd143;
#400 gamma=32'd5;row=32'd486;
#400 gamma=32'd2;row=32'd198;
#400 gamma=32'd1;row=32'd536;
#400 gamma=32'd3;row=32'd411;
#400 gamma=32'd1;row=32'd232;
#400 gamma=32'd5;row=32'd238;
#400 gamma=32'd5;row=32'd374;
#400 gamma=32'd4;row=32'd168;
#400 gamma=32'd4;row=32'd55;
#400 gamma=32'd2;row=32'd107;
#400 gamma=32'd3;row=32'd389;
#400 gamma=32'd2;row=32'd252;
#400 gamma=32'd1;row=32'd430;
#400 gamma=32'd2;row=32'd181;
#400 gamma=32'd3;row=32'd426;
#400 gamma=32'd5;row=32'd29;
#400 gamma=32'd5;row=32'd56;
#400 gamma=32'd1;row=32'd28;
#400 gamma=32'd1;row=32'd472;
#400 gamma=32'd5;row=32'd324;
#400 gamma=32'd2;row=32'd151;
#400 gamma=32'd3;row=32'd243;
#400 gamma=32'd1;row=32'd417;
#400 gamma=32'd3;row=32'd172;
#400 gamma=32'd3;row=32'd123;
#400 gamma=32'd1;row=32'd126;
#400 gamma=32'd1;row=32'd398;
#400 gamma=32'd1;row=32'd71;
#400 gamma=32'd3;row=32'd335;
#400 gamma=32'd2;row=32'd192;
#400 gamma=32'd2;row=32'd401;
#400 gamma=32'd1;row=32'd512;
#400 gamma=32'd1;row=32'd10;
#400 gamma=32'd3;row=32'd357;
#400 gamma=32'd2;row=32'd467;
#400 gamma=32'd5;row=32'd355;
#400 gamma=32'd5;row=32'd339;
#400 gamma=32'd1;row=32'd54;
#400 gamma=32'd2;row=32'd474;
#400 gamma=32'd1;row=32'd356;
#400 gamma=32'd2;row=32'd123;
#400 gamma=32'd5;row=32'd505;
#400 gamma=32'd3;row=32'd386;
#400 gamma=32'd1;row=32'd128;
#400 gamma=32'd2;row=32'd285;
#400 gamma=32'd3;row=32'd171;
#400 gamma=32'd5;row=32'd263;
#400 gamma=32'd2;row=32'd62;
#400 gamma=32'd4;row=32'd58;
#400 gamma=32'd2;row=32'd508;
#400 gamma=32'd2;row=32'd323;
#400 gamma=32'd4;row=32'd386;
#400 gamma=32'd4;row=32'd394;
#400 gamma=32'd4;row=32'd483;
#400 gamma=32'd2;row=32'd152;
#400 gamma=32'd4;row=32'd169;
#400 gamma=32'd5;row=32'd215;
#400 gamma=32'd3;row=32'd416;
#400 gamma=32'd3;row=32'd447;
#400 gamma=32'd5;row=32'd90;
#400 gamma=32'd2;row=32'd541;
#400 gamma=32'd4;row=32'd0;
#400 gamma=32'd4;row=32'd323;
#400 gamma=32'd2;row=32'd13;
#400 gamma=32'd3;row=32'd553;
#400 gamma=32'd2;row=32'd359;
#400 gamma=32'd1;row=32'd403;
#400 gamma=32'd1;row=32'd466;
#400 gamma=32'd4;row=32'd178;
#400 gamma=32'd4;row=32'd208;
#400 gamma=32'd2;row=32'd112;
#400 gamma=32'd3;row=32'd137;
#400 gamma=32'd2;row=32'd532;
#400 gamma=32'd1;row=32'd206;
#400 gamma=32'd4;row=32'd436;
#400 gamma=32'd4;row=32'd189;
#400 gamma=32'd5;row=32'd166;
#400 gamma=32'd5;row=32'd183;
#400 gamma=32'd4;row=32'd239;
#400 gamma=32'd5;row=32'd21;
#400 gamma=32'd4;row=32'd327;
#400 gamma=32'd4;row=32'd20;
#400 gamma=32'd5;row=32'd187;
#400 gamma=32'd4;row=32'd362;
#400 gamma=32'd5;row=32'd446;
#400 gamma=32'd5;row=32'd235;
#400 gamma=32'd2;row=32'd343;
#400 gamma=32'd5;row=32'd47;
#400 gamma=32'd5;row=32'd121;
#400 gamma=32'd2;row=32'd344;
#400 gamma=32'd3;row=32'd249;
#400 gamma=32'd2;row=32'd552;
#400 gamma=32'd2;row=32'd25;
#400 gamma=32'd1;row=32'd287;
#400 gamma=32'd2;row=32'd331;
#400 gamma=32'd3;row=32'd155;
#400 gamma=32'd4;row=32'd2;
#400 gamma=32'd2;row=32'd542;
#400 gamma=32'd4;row=32'd506;
#400 gamma=32'd2;row=32'd458;
#400 gamma=32'd1;row=32'd28;
#400 gamma=32'd2;row=32'd451;
#400 gamma=32'd1;row=32'd255;
#400 gamma=32'd4;row=32'd417;
#400 gamma=32'd3;row=32'd84;
#400 gamma=32'd1;row=32'd165;
#400 gamma=32'd3;row=32'd205;
#400 gamma=32'd3;row=32'd403;
#400 gamma=32'd2;row=32'd355;
#400 gamma=32'd3;row=32'd403;
#400 gamma=32'd5;row=32'd17;
#400 gamma=32'd3;row=32'd56;
#400 gamma=32'd3;row=32'd373;
#400 gamma=32'd1;row=32'd46;
#400 gamma=32'd1;row=32'd67;
#400 gamma=32'd2;row=32'd376;
#400 gamma=32'd2;row=32'd153;
#400 gamma=32'd4;row=32'd206;
#400 gamma=32'd5;row=32'd489;
#400 gamma=32'd5;row=32'd57;
#400 gamma=32'd3;row=32'd33;
#400 gamma=32'd1;row=32'd121;
#400 gamma=32'd2;row=32'd370;
#400 gamma=32'd2;row=32'd300;
#400 gamma=32'd2;row=32'd36;
#400 gamma=32'd1;row=32'd73;
#400 gamma=32'd3;row=32'd117;
#400 gamma=32'd3;row=32'd97;
#400 gamma=32'd3;row=32'd98;
#400 gamma=32'd2;row=32'd370;
#400 gamma=32'd3;row=32'd223;
#400 gamma=32'd5;row=32'd224;
#400 gamma=32'd5;row=32'd133;
#400 gamma=32'd1;row=32'd430;
#400 gamma=32'd1;row=32'd325;
#400 gamma=32'd2;row=32'd340;
#400 gamma=32'd3;row=32'd91;
#400 gamma=32'd3;row=32'd52;
#400 gamma=32'd1;row=32'd361;
#400 gamma=32'd5;row=32'd507;
#400 gamma=32'd2;row=32'd91;
#400 gamma=32'd4;row=32'd167;
#400 gamma=32'd1;row=32'd268;
#400 gamma=32'd1;row=32'd157;
#400 gamma=32'd4;row=32'd244;
#400 gamma=32'd1;row=32'd198;
#400 gamma=32'd2;row=32'd30;
#400 gamma=32'd4;row=32'd138;
#400 gamma=32'd5;row=32'd1;
#400 gamma=32'd4;row=32'd249;
#400 gamma=32'd3;row=32'd172;
#400 gamma=32'd2;row=32'd271;
#400 gamma=32'd5;row=32'd428;
#400 gamma=32'd2;row=32'd87;
#400 gamma=32'd5;row=32'd118;
#400 gamma=32'd2;row=32'd508;
#400 gamma=32'd1;row=32'd26;
#400 gamma=32'd4;row=32'd254;
#400 gamma=32'd1;row=32'd489;
#400 gamma=32'd1;row=32'd534;
#400 gamma=32'd2;row=32'd433;
#400 gamma=32'd5;row=32'd37;
#400 gamma=32'd2;row=32'd79;
#400 gamma=32'd3;row=32'd168;
#400 gamma=32'd5;row=32'd1;
#400 gamma=32'd5;row=32'd94;
#400 gamma=32'd2;row=32'd312;
#400 gamma=32'd3;row=32'd395;
#400 gamma=32'd2;row=32'd489;
#400 gamma=32'd1;row=32'd58;
#400 gamma=32'd1;row=32'd435;
#400 gamma=32'd3;row=32'd131;
#400 gamma=32'd3;row=32'd80;
#400 gamma=32'd3;row=32'd64;
#400 gamma=32'd5;row=32'd251;
#400 gamma=32'd5;row=32'd328;
#400 gamma=32'd1;row=32'd96;
#400 gamma=32'd3;row=32'd89;
#400 gamma=32'd4;row=32'd468;
#400 gamma=32'd4;row=32'd385;
#400 gamma=32'd2;row=32'd451;
#400 gamma=32'd2;row=32'd196;
#400 gamma=32'd5;row=32'd533;
#400 gamma=32'd2;row=32'd311;
#400 gamma=32'd4;row=32'd412;
#400 gamma=32'd1;row=32'd93;
#400 gamma=32'd2;row=32'd434;
#400 gamma=32'd3;row=32'd234;
#400 gamma=32'd1;row=32'd189;
#400 gamma=32'd2;row=32'd456;
#400 gamma=32'd3;row=32'd101;
#400 gamma=32'd2;row=32'd424;
#400 gamma=32'd1;row=32'd32;
#400 gamma=32'd3;row=32'd186;
#400 gamma=32'd1;row=32'd386;
#400 gamma=32'd2;row=32'd426;
#400 gamma=32'd1;row=32'd82;
#400 gamma=32'd4;row=32'd261;
#400 gamma=32'd4;row=32'd330;
#400 gamma=32'd3;row=32'd165;
#400 gamma=32'd3;row=32'd390;
#400 gamma=32'd1;row=32'd204;
#400 gamma=32'd4;row=32'd201;
#400 gamma=32'd2;row=32'd229;
#400 gamma=32'd2;row=32'd37;
#400 gamma=32'd5;row=32'd132;
#400 gamma=32'd2;row=32'd420;
#400 gamma=32'd2;row=32'd20;
#400 gamma=32'd2;row=32'd274;
#400 gamma=32'd3;row=32'd330;
#400 gamma=32'd4;row=32'd324;
#400 gamma=32'd4;row=32'd2;
#400 gamma=32'd2;row=32'd408;
#400 gamma=32'd3;row=32'd447;
#400 gamma=32'd4;row=32'd359;
#400 gamma=32'd2;row=32'd335;
#400 gamma=32'd3;row=32'd22;
#400 gamma=32'd2;row=32'd154;
#400 gamma=32'd5;row=32'd168;
#400 gamma=32'd2;row=32'd231;
#400 gamma=32'd3;row=32'd257;
#400 gamma=32'd3;row=32'd494;
#400 gamma=32'd5;row=32'd476;
#400 gamma=32'd2;row=32'd218;
#400 gamma=32'd4;row=32'd372;
#400 gamma=32'd1;row=32'd11;
#400 gamma=32'd5;row=32'd510;
#400 gamma=32'd5;row=32'd36;
#400 gamma=32'd2;row=32'd431;
#400 gamma=32'd5;row=32'd128;
#400 gamma=32'd4;row=32'd284;
#400 gamma=32'd2;row=32'd319;
#400 gamma=32'd1;row=32'd436;
#400 gamma=32'd1;row=32'd373;
#400 gamma=32'd5;row=32'd88;
#400 gamma=32'd1;row=32'd219;
#400 gamma=32'd5;row=32'd319;
#400 gamma=32'd4;row=32'd180;
#400 gamma=32'd1;row=32'd244;
#400 gamma=32'd4;row=32'd467;
#400 gamma=32'd3;row=32'd478;
#400 gamma=32'd4;row=32'd324;
#400 gamma=32'd3;row=32'd386;
#400 gamma=32'd3;row=32'd256;
#400 gamma=32'd3;row=32'd418;
#400 gamma=32'd4;row=32'd455;
#400 gamma=32'd1;row=32'd323;
#400 gamma=32'd5;row=32'd140;
#400 gamma=32'd4;row=32'd322;
#400 gamma=32'd1;row=32'd550;
#400 gamma=32'd5;row=32'd242;
#400 gamma=32'd5;row=32'd18;
#400 gamma=32'd5;row=32'd139;
#400 gamma=32'd2;row=32'd422;
#400 gamma=32'd5;row=32'd107;
#400 gamma=32'd2;row=32'd451;
#400 gamma=32'd5;row=32'd72;
#400 gamma=32'd4;row=32'd477;
#400 gamma=32'd3;row=32'd487;
#400 gamma=32'd2;row=32'd296;
#400 gamma=32'd1;row=32'd71;
#400 gamma=32'd3;row=32'd187;
#400 gamma=32'd4;row=32'd69;
#400 gamma=32'd2;row=32'd156;
#400 gamma=32'd3;row=32'd512;
#400 gamma=32'd5;row=32'd386;
#400 gamma=32'd3;row=32'd455;
#400 gamma=32'd3;row=32'd98;
#400 gamma=32'd5;row=32'd24;
#400 gamma=32'd4;row=32'd246;
#400 gamma=32'd1;row=32'd495;
#400 gamma=32'd5;row=32'd500;
#400 gamma=32'd4;row=32'd554;
#400 gamma=32'd1;row=32'd91;
#400 gamma=32'd1;row=32'd294;
#400 gamma=32'd4;row=32'd541;
#400 gamma=32'd5;row=32'd62;
#400 gamma=32'd4;row=32'd374;
#400 gamma=32'd3;row=32'd549;
#400 gamma=32'd1;row=32'd249;
#400 gamma=32'd1;row=32'd454;
#400 gamma=32'd2;row=32'd310;
#400 gamma=32'd5;row=32'd452;
#400 gamma=32'd3;row=32'd109;
#400 gamma=32'd2;row=32'd138;
#400 gamma=32'd2;row=32'd145;
#400 gamma=32'd4;row=32'd319;
#400 gamma=32'd1;row=32'd36;
#400 gamma=32'd2;row=32'd319;
#400 gamma=32'd1;row=32'd230;
#400 gamma=32'd2;row=32'd367;
#400 gamma=32'd5;row=32'd37;
#400 gamma=32'd5;row=32'd408;
#400 gamma=32'd2;row=32'd535;
#400 gamma=32'd3;row=32'd248;
#400 gamma=32'd2;row=32'd432;
#400 gamma=32'd3;row=32'd244;
#400 gamma=32'd4;row=32'd417;
#400 gamma=32'd2;row=32'd258;
#400 gamma=32'd4;row=32'd141;
#400 gamma=32'd5;row=32'd225;
#400 gamma=32'd3;row=32'd470;
#400 gamma=32'd3;row=32'd212;
#400 gamma=32'd3;row=32'd418;
#400 gamma=32'd3;row=32'd383;
#400 gamma=32'd5;row=32'd390;
#400 gamma=32'd3;row=32'd136;
#400 gamma=32'd1;row=32'd121;
#400 gamma=32'd2;row=32'd498;
#400 gamma=32'd2;row=32'd98;
#400 gamma=32'd1;row=32'd337;
#400 gamma=32'd1;row=32'd340;
#400 gamma=32'd5;row=32'd91;
#400 gamma=32'd4;row=32'd232;
#400 gamma=32'd3;row=32'd250;
#400 gamma=32'd2;row=32'd438;
#400 gamma=32'd1;row=32'd237;
#400 gamma=32'd1;row=32'd200;
#400 gamma=32'd2;row=32'd234;
#400 gamma=32'd5;row=32'd468;
#400 gamma=32'd5;row=32'd0;
#400 gamma=32'd5;row=32'd108;
#400 gamma=32'd3;row=32'd283;
#400 gamma=32'd2;row=32'd170;
#400 gamma=32'd2;row=32'd16;
#400 gamma=32'd3;row=32'd64;
#400 gamma=32'd4;row=32'd111;
#400 gamma=32'd1;row=32'd411;
#400 gamma=32'd5;row=32'd550;
#400 gamma=32'd3;row=32'd338;
#400 gamma=32'd3;row=32'd349;
#400 gamma=32'd5;row=32'd299;
#400 gamma=32'd3;row=32'd418;
#400 gamma=32'd2;row=32'd50;
#400 gamma=32'd1;row=32'd555;
#400 gamma=32'd5;row=32'd130;
#400 gamma=32'd1;row=32'd165;
#400 gamma=32'd3;row=32'd314;
#400 gamma=32'd2;row=32'd136;
#400 gamma=32'd1;row=32'd154;
#400 gamma=32'd2;row=32'd102;
#400 gamma=32'd4;row=32'd158;
#400 gamma=32'd3;row=32'd541;
#400 gamma=32'd5;row=32'd218;
#400 gamma=32'd4;row=32'd142;
#400 gamma=32'd5;row=32'd354;
#400 gamma=32'd3;row=32'd505;
#400 gamma=32'd2;row=32'd126;
#400 gamma=32'd3;row=32'd148;
#400 gamma=32'd1;row=32'd466;
#400 gamma=32'd4;row=32'd142;
#400 gamma=32'd4;row=32'd51;
#400 gamma=32'd4;row=32'd465;
#400 gamma=32'd1;row=32'd78;
#400 gamma=32'd5;row=32'd334;
#400 gamma=32'd2;row=32'd47;
#400 gamma=32'd1;row=32'd335;
#400 gamma=32'd5;row=32'd90;
#400 gamma=32'd5;row=32'd215;
#400 gamma=32'd4;row=32'd82;
#400 gamma=32'd5;row=32'd373;
#400 gamma=32'd2;row=32'd56;
#400 gamma=32'd2;row=32'd91;
#400 gamma=32'd4;row=32'd352;
#400 gamma=32'd4;row=32'd557;
#400 gamma=32'd1;row=32'd197;
#400 gamma=32'd1;row=32'd26;
#400 gamma=32'd1;row=32'd546;
#400 gamma=32'd4;row=32'd321;
#400 gamma=32'd2;row=32'd92;
#400 gamma=32'd2;row=32'd181;
#400 gamma=32'd3;row=32'd456;
#400 gamma=32'd3;row=32'd301;
#400 gamma=32'd2;row=32'd196;
#400 gamma=32'd3;row=32'd359;
#400 gamma=32'd3;row=32'd328;
#400 gamma=32'd1;row=32'd483;
#400 gamma=32'd1;row=32'd261;
#400 gamma=32'd1;row=32'd241;
#400 gamma=32'd1;row=32'd38;
#400 gamma=32'd1;row=32'd237;
#400 gamma=32'd1;row=32'd65;
#400 gamma=32'd4;row=32'd40;
#400 gamma=32'd4;row=32'd26;
#400 gamma=32'd5;row=32'd454;
#400 gamma=32'd2;row=32'd43;
#400 gamma=32'd4;row=32'd552;
#400 gamma=32'd1;row=32'd501;
#400 gamma=32'd5;row=32'd143;
#400 gamma=32'd5;row=32'd145;
#400 gamma=32'd5;row=32'd52;
#400 gamma=32'd4;row=32'd212;
#400 gamma=32'd1;row=32'd60;
#400 gamma=32'd1;row=32'd154;
#400 gamma=32'd3;row=32'd153;
#400 gamma=32'd5;row=32'd231;
#400 gamma=32'd3;row=32'd75;
#400 gamma=32'd1;row=32'd68;
#400 gamma=32'd1;row=32'd313;
#400 gamma=32'd3;row=32'd468;
#400 gamma=32'd5;row=32'd548;
#400 gamma=32'd4;row=32'd491;
#400 gamma=32'd1;row=32'd343;
#400 gamma=32'd4;row=32'd98;
#400 gamma=32'd4;row=32'd30;
#400 gamma=32'd5;row=32'd465;
#400 gamma=32'd4;row=32'd306;
#400 gamma=32'd4;row=32'd426;
#400 gamma=32'd3;row=32'd466;
#400 gamma=32'd3;row=32'd488;
#400 gamma=32'd3;row=32'd223;
#400 gamma=32'd4;row=32'd449;
#400 gamma=32'd5;row=32'd431;
#400 gamma=32'd1;row=32'd382;
#400 gamma=32'd1;row=32'd412;
#400 gamma=32'd3;row=32'd168;
#400 gamma=32'd3;row=32'd177;
#400 gamma=32'd4;row=32'd527;
#400 gamma=32'd5;row=32'd167;
#400 gamma=32'd5;row=32'd93;
#400 gamma=32'd1;row=32'd366;
#400 gamma=32'd2;row=32'd168;
#400 gamma=32'd3;row=32'd13;
#400 gamma=32'd1;row=32'd242;
#400 gamma=32'd3;row=32'd9;
#400 gamma=32'd4;row=32'd520;
#400 gamma=32'd3;row=32'd31;
#400 gamma=32'd5;row=32'd47;
#400 gamma=32'd1;row=32'd105;
#400 gamma=32'd3;row=32'd498;
#400 gamma=32'd2;row=32'd36;
#400 gamma=32'd1;row=32'd386;
#400 gamma=32'd3;row=32'd196;
#400 gamma=32'd5;row=32'd269;
#400 gamma=32'd3;row=32'd308;
#400 gamma=32'd1;row=32'd98;
#400 gamma=32'd5;row=32'd399;
#400 gamma=32'd4;row=32'd544;
#400 gamma=32'd4;row=32'd93;
#400 gamma=32'd5;row=32'd478;
#400 gamma=32'd1;row=32'd385;
#400 gamma=32'd1;row=32'd476;
#400 gamma=32'd1;row=32'd96;
#400 gamma=32'd2;row=32'd234;
#400 gamma=32'd4;row=32'd414;
#400 gamma=32'd4;row=32'd481;
#400 gamma=32'd3;row=32'd493;
#400 gamma=32'd1;row=32'd129;
#400 gamma=32'd3;row=32'd554;
#400 gamma=32'd5;row=32'd3;
#400 gamma=32'd5;row=32'd378;
#400 gamma=32'd1;row=32'd287;
#400 gamma=32'd4;row=32'd282;
#400 gamma=32'd3;row=32'd270;
#400 gamma=32'd2;row=32'd544;
#400 gamma=32'd4;row=32'd152;
#400 gamma=32'd1;row=32'd175;
#400 gamma=32'd1;row=32'd104;
#400 gamma=32'd3;row=32'd431;
#400 gamma=32'd2;row=32'd509;
#400 gamma=32'd1;row=32'd180;
#400 gamma=32'd2;row=32'd86;
#400 gamma=32'd3;row=32'd35;
#400 gamma=32'd2;row=32'd295;
#400 gamma=32'd1;row=32'd223;
#400 gamma=32'd5;row=32'd94;
#400 gamma=32'd5;row=32'd503;
#400 gamma=32'd3;row=32'd382;
#400 gamma=32'd3;row=32'd368;
#400 gamma=32'd2;row=32'd528;
#400 gamma=32'd1;row=32'd15;
#400 gamma=32'd5;row=32'd101;
#400 gamma=32'd2;row=32'd120;
#400 gamma=32'd3;row=32'd469;
#400 gamma=32'd2;row=32'd556;
#400 gamma=32'd3;row=32'd171;
#400 gamma=32'd4;row=32'd328;
#400 gamma=32'd2;row=32'd150;
#400 gamma=32'd2;row=32'd226;
#400 gamma=32'd2;row=32'd22;
#400 gamma=32'd5;row=32'd85;
#400 gamma=32'd4;row=32'd117;
#400 gamma=32'd2;row=32'd468;
#400 gamma=32'd3;row=32'd491;
#400 gamma=32'd4;row=32'd544;
#400 gamma=32'd5;row=32'd402;
#400 gamma=32'd2;row=32'd500;
#400 gamma=32'd5;row=32'd113;
#400 gamma=32'd5;row=32'd24;
#400 gamma=32'd3;row=32'd502;
#400 gamma=32'd1;row=32'd405;
#400 gamma=32'd4;row=32'd265;
#400 gamma=32'd5;row=32'd177;
#400 gamma=32'd3;row=32'd217;
#400 gamma=32'd1;row=32'd164;
#400 gamma=32'd3;row=32'd85;
#400 gamma=32'd2;row=32'd120;
#400 gamma=32'd2;row=32'd457;
#400 gamma=32'd2;row=32'd172;
#400 gamma=32'd1;row=32'd293;
#400 gamma=32'd1;row=32'd294;
#400 gamma=32'd5;row=32'd216;
#400 gamma=32'd1;row=32'd435;
#400 gamma=32'd4;row=32'd434;
#400 gamma=32'd3;row=32'd487;
#400 gamma=32'd3;row=32'd553;
#400 gamma=32'd3;row=32'd48;
#400 gamma=32'd3;row=32'd403;
#400 gamma=32'd4;row=32'd62;
#400 gamma=32'd4;row=32'd84;
#400 gamma=32'd3;row=32'd62;
#400 gamma=32'd3;row=32'd218;
#400 gamma=32'd2;row=32'd118;
#400 gamma=32'd3;row=32'd154;
#400 gamma=32'd2;row=32'd442;
#400 gamma=32'd5;row=32'd268;
#400 gamma=32'd2;row=32'd558;
#400 gamma=32'd1;row=32'd42;
#400 gamma=32'd2;row=32'd112;
#400 gamma=32'd4;row=32'd487;
#400 gamma=32'd2;row=32'd328;
#400 gamma=32'd1;row=32'd180;
#400 gamma=32'd2;row=32'd376;
#400 gamma=32'd5;row=32'd81;
#400 gamma=32'd3;row=32'd108;
#400 gamma=32'd1;row=32'd256;
#400 gamma=32'd5;row=32'd472;
#400 gamma=32'd5;row=32'd212;
#400 gamma=32'd5;row=32'd325;
#400 gamma=32'd2;row=32'd522;
#400 gamma=32'd1;row=32'd402;
#400 gamma=32'd1;row=32'd341;
#400 gamma=32'd4;row=32'd133;
#400 gamma=32'd4;row=32'd415;
#400 gamma=32'd4;row=32'd230;
#400 gamma=32'd1;row=32'd44;
#400 gamma=32'd2;row=32'd207;
#400 gamma=32'd4;row=32'd103;
#400 gamma=32'd2;row=32'd381;
#400 gamma=32'd1;row=32'd9;
#400 gamma=32'd5;row=32'd213;
#400 gamma=32'd3;row=32'd499;
#400 gamma=32'd1;row=32'd303;
#400 gamma=32'd4;row=32'd86;
#400 gamma=32'd4;row=32'd196;
#400 gamma=32'd5;row=32'd527;
#400 gamma=32'd1;row=32'd357;
#400 gamma=32'd2;row=32'd355;
#400 gamma=32'd5;row=32'd374;
#400 gamma=32'd4;row=32'd54;
#400 gamma=32'd3;row=32'd32;
#400 gamma=32'd4;row=32'd422;
#400 gamma=32'd1;row=32'd276;
#400 gamma=32'd1;row=32'd474;
#400 gamma=32'd5;row=32'd325;
#400 gamma=32'd2;row=32'd192;
#400 gamma=32'd3;row=32'd372;
#400 gamma=32'd4;row=32'd435;
#400 gamma=32'd5;row=32'd489;
#400 gamma=32'd5;row=32'd395;
#400 gamma=32'd3;row=32'd495;
#400 gamma=32'd4;row=32'd395;
#400 gamma=32'd2;row=32'd7;
#400 gamma=32'd1;row=32'd259;
#400 gamma=32'd4;row=32'd29;
#400 gamma=32'd3;row=32'd63;
#400 gamma=32'd3;row=32'd238;
#400 gamma=32'd2;row=32'd500;
#400 gamma=32'd5;row=32'd90;
#400 gamma=32'd5;row=32'd18;
#400 gamma=32'd5;row=32'd320;
#400 gamma=32'd5;row=32'd445;
#400 gamma=32'd3;row=32'd181;
#400 gamma=32'd2;row=32'd531;
#400 gamma=32'd2;row=32'd495;
#400 gamma=32'd5;row=32'd61;
#400 gamma=32'd3;row=32'd316;
#400 gamma=32'd3;row=32'd356;
#400 gamma=32'd2;row=32'd554;
#400 gamma=32'd3;row=32'd156;
#400 gamma=32'd5;row=32'd552;
#400 gamma=32'd4;row=32'd160;
#400 gamma=32'd1;row=32'd348;
#400 gamma=32'd2;row=32'd121;
#400 gamma=32'd5;row=32'd460;
#400 gamma=32'd3;row=32'd157;
#400 gamma=32'd5;row=32'd330;
#400 gamma=32'd4;row=32'd82;
#400 gamma=32'd2;row=32'd22;
#400 gamma=32'd2;row=32'd210;
#400 gamma=32'd4;row=32'd480;
#400 gamma=32'd5;row=32'd433;
#400 gamma=32'd5;row=32'd421;
#400 gamma=32'd2;row=32'd19;
#400 gamma=32'd1;row=32'd237;
#400 gamma=32'd4;row=32'd265;
#400 gamma=32'd1;row=32'd508;
#400 gamma=32'd4;row=32'd441;
#400 gamma=32'd4;row=32'd122;
#400 gamma=32'd5;row=32'd45;
#400 gamma=32'd4;row=32'd428;
#400 gamma=32'd2;row=32'd239;
#400 gamma=32'd4;row=32'd93;
#400 gamma=32'd5;row=32'd318;
#400 gamma=32'd2;row=32'd164;
#400 gamma=32'd2;row=32'd222;
#400 gamma=32'd1;row=32'd83;
#400 gamma=32'd3;row=32'd357;
#400 gamma=32'd3;row=32'd500;
#400 gamma=32'd3;row=32'd84;
#400 gamma=32'd1;row=32'd22;
#400 gamma=32'd3;row=32'd536;
#400 gamma=32'd2;row=32'd100;
#400 gamma=32'd4;row=32'd278;
#400 gamma=32'd2;row=32'd170;
#400 gamma=32'd4;row=32'd312;
#400 gamma=32'd5;row=32'd62;
#400 gamma=32'd5;row=32'd13;
#400 gamma=32'd4;row=32'd79;
#400 gamma=32'd1;row=32'd403;
#400 gamma=32'd5;row=32'd479;
#400 gamma=32'd1;row=32'd423;
#400 gamma=32'd4;row=32'd287;
#400 gamma=32'd3;row=32'd488;
#400 gamma=32'd1;row=32'd383;
#400 gamma=32'd1;row=32'd185;
#400 gamma=32'd1;row=32'd94;
#400 gamma=32'd5;row=32'd332;
#400 gamma=32'd3;row=32'd499;
#400 gamma=32'd4;row=32'd530;
#400 gamma=32'd1;row=32'd498;
#400 gamma=32'd2;row=32'd38;
#400 gamma=32'd1;row=32'd547;
#400 gamma=32'd2;row=32'd455;
#400 gamma=32'd4;row=32'd101;
#400 gamma=32'd3;row=32'd108;
#400 gamma=32'd2;row=32'd26;
#400 gamma=32'd1;row=32'd355;
#400 gamma=32'd4;row=32'd272;
#400 gamma=32'd4;row=32'd405;
#400 gamma=32'd4;row=32'd322;
#400 gamma=32'd4;row=32'd145;
#400 gamma=32'd2;row=32'd258;
#400 gamma=32'd4;row=32'd256;
#400 gamma=32'd4;row=32'd157;
#400 gamma=32'd3;row=32'd196;
#400 gamma=32'd5;row=32'd127;
#400 gamma=32'd4;row=32'd0;
#400 gamma=32'd5;row=32'd537;
#400 gamma=32'd4;row=32'd510;
#400 gamma=32'd5;row=32'd328;
#400 gamma=32'd4;row=32'd151;
#400 gamma=32'd2;row=32'd242;
#400 gamma=32'd2;row=32'd152;
#400 gamma=32'd1;row=32'd478;
#400 gamma=32'd2;row=32'd263;
#400 gamma=32'd5;row=32'd221;
#400 gamma=32'd3;row=32'd454;
#400 gamma=32'd1;row=32'd2;
#400 gamma=32'd5;row=32'd295;
#400 gamma=32'd1;row=32'd439;
#400 gamma=32'd2;row=32'd536;
#400 gamma=32'd1;row=32'd424;
#400 gamma=32'd5;row=32'd89;
#400 gamma=32'd2;row=32'd427;
#400 gamma=32'd4;row=32'd143;
#400 gamma=32'd2;row=32'd317;
#400 gamma=32'd1;row=32'd378;
#400 gamma=32'd1;row=32'd438;
#400 gamma=32'd4;row=32'd442;
#400 gamma=32'd4;row=32'd243;
#400 gamma=32'd4;row=32'd76;
#400 gamma=32'd3;row=32'd392;
#400 gamma=32'd1;row=32'd143;
#400 gamma=32'd2;row=32'd342;
#400 gamma=32'd2;row=32'd132;
#400 gamma=32'd3;row=32'd295;
#400 gamma=32'd3;row=32'd494;
#400 gamma=32'd1;row=32'd430;
#400 gamma=32'd4;row=32'd379;
#400 gamma=32'd5;row=32'd10;
#400 gamma=32'd3;row=32'd541;
#400 gamma=32'd5;row=32'd287;
#400 gamma=32'd4;row=32'd116;
#400 gamma=32'd3;row=32'd131;
#400 gamma=32'd1;row=32'd14;
#400 gamma=32'd1;row=32'd528;
#400 gamma=32'd5;row=32'd277;
#400 gamma=32'd2;row=32'd125;
#400 gamma=32'd5;row=32'd198;
#400 gamma=32'd1;row=32'd55;
#400 gamma=32'd5;row=32'd68;
#400 gamma=32'd3;row=32'd5;
#400 gamma=32'd2;row=32'd317;
#400 gamma=32'd4;row=32'd21;
#400 gamma=32'd2;row=32'd554;
#400 gamma=32'd1;row=32'd383;
#400 gamma=32'd4;row=32'd525;
#400 gamma=32'd2;row=32'd484;
#400 gamma=32'd3;row=32'd212;
#400 gamma=32'd2;row=32'd374;
#400 gamma=32'd2;row=32'd412;
#400 gamma=32'd4;row=32'd211;
#400 gamma=32'd4;row=32'd78;
#400 gamma=32'd3;row=32'd359;
#400 gamma=32'd4;row=32'd3;
#400 gamma=32'd4;row=32'd167;
#400 gamma=32'd4;row=32'd327;
#400 gamma=32'd4;row=32'd35;
#400 gamma=32'd1;row=32'd245;
#400 gamma=32'd5;row=32'd56;
#400 gamma=32'd3;row=32'd514;
#400 gamma=32'd1;row=32'd479;
#400 gamma=32'd3;row=32'd517;
#400 gamma=32'd3;row=32'd326;
#400 gamma=32'd2;row=32'd126;
#400 gamma=32'd4;row=32'd152;
#400 gamma=32'd4;row=32'd328;
#400 gamma=32'd1;row=32'd284;
#400 gamma=32'd2;row=32'd229;
#400 gamma=32'd5;row=32'd559;
#400 gamma=32'd1;row=32'd7;
#400 gamma=32'd3;row=32'd52;
#400 gamma=32'd4;row=32'd21;
#400 gamma=32'd3;row=32'd228;
#400 gamma=32'd1;row=32'd319;
#400 gamma=32'd5;row=32'd516;
#400 gamma=32'd1;row=32'd414;
#400 gamma=32'd3;row=32'd205;
#400 gamma=32'd1;row=32'd275;
#400 gamma=32'd5;row=32'd5;
#400 gamma=32'd3;row=32'd388;
#400 gamma=32'd2;row=32'd546;
#400 gamma=32'd5;row=32'd284;
#400 gamma=32'd2;row=32'd223;
#400 gamma=32'd2;row=32'd230;
#400 gamma=32'd5;row=32'd409;
#400 gamma=32'd5;row=32'd299;
#400 gamma=32'd3;row=32'd182;
#400 gamma=32'd2;row=32'd211;
#400 gamma=32'd4;row=32'd307;
#400 gamma=32'd5;row=32'd315;
#400 gamma=32'd5;row=32'd256;
#400 gamma=32'd5;row=32'd268;
#400 gamma=32'd3;row=32'd277;
#400 gamma=32'd3;row=32'd465;
#400 gamma=32'd5;row=32'd243;
#400 gamma=32'd3;row=32'd334;
#400 gamma=32'd2;row=32'd510;
#400 gamma=32'd3;row=32'd289;
#400 gamma=32'd1;row=32'd96;
#400 gamma=32'd1;row=32'd463;
#400 gamma=32'd4;row=32'd101;
#400 gamma=32'd5;row=32'd492;
#400 gamma=32'd1;row=32'd349;
#400 gamma=32'd2;row=32'd73;
#400 gamma=32'd4;row=32'd383;
#400 gamma=32'd4;row=32'd160;
#400 gamma=32'd4;row=32'd513;
#400 gamma=32'd3;row=32'd210;
#400 gamma=32'd2;row=32'd548;
#400 gamma=32'd2;row=32'd321;
#400 gamma=32'd3;row=32'd302;
#400 gamma=32'd5;row=32'd136;
#400 gamma=32'd3;row=32'd384;
#400 gamma=32'd2;row=32'd104;
#400 gamma=32'd5;row=32'd11;
#400 gamma=32'd4;row=32'd478;
#400 gamma=32'd1;row=32'd244;
#400 gamma=32'd2;row=32'd212;
#400 gamma=32'd5;row=32'd496;
#400 gamma=32'd1;row=32'd417;
#400 gamma=32'd2;row=32'd360;
#400 gamma=32'd3;row=32'd338;
#400 gamma=32'd1;row=32'd317;
#400 gamma=32'd3;row=32'd31;
#400 gamma=32'd3;row=32'd46;
#400 gamma=32'd3;row=32'd60;
#400 gamma=32'd2;row=32'd56;
#400 gamma=32'd1;row=32'd315;
#400 gamma=32'd3;row=32'd376;
#400 gamma=32'd5;row=32'd10;
#400 gamma=32'd2;row=32'd465;
#400 gamma=32'd3;row=32'd167;
#400 gamma=32'd2;row=32'd358;
#400 gamma=32'd2;row=32'd310;
#400 gamma=32'd4;row=32'd240;
#400 gamma=32'd1;row=32'd364;
#400 gamma=32'd3;row=32'd554;
#400 gamma=32'd5;row=32'd81;
#400 gamma=32'd5;row=32'd231;
#400 gamma=32'd5;row=32'd6;
#400 gamma=32'd2;row=32'd402;
#400 gamma=32'd1;row=32'd200;
#400 gamma=32'd2;row=32'd511;
#400 gamma=32'd5;row=32'd471;
#400 gamma=32'd3;row=32'd75;
#400 gamma=32'd4;row=32'd349;
#400 gamma=32'd5;row=32'd165;
#400 gamma=32'd3;row=32'd457;
#400 gamma=32'd5;row=32'd151;
#400 gamma=32'd4;row=32'd74;
#400 gamma=32'd5;row=32'd4;
#400 gamma=32'd3;row=32'd266;
#400 gamma=32'd3;row=32'd186;
#400 gamma=32'd5;row=32'd314;
#400 gamma=32'd1;row=32'd359;
#400 gamma=32'd4;row=32'd139;
#400 gamma=32'd1;row=32'd370;
#400 gamma=32'd1;row=32'd231;
#400 gamma=32'd1;row=32'd473;
#400 gamma=32'd3;row=32'd122;
#400 gamma=32'd4;row=32'd529;
#400 gamma=32'd5;row=32'd223;
#400 gamma=32'd5;row=32'd540;
#400 gamma=32'd1;row=32'd277;
#400 gamma=32'd4;row=32'd46;
#400 gamma=32'd2;row=32'd155;
#400 gamma=32'd4;row=32'd399;
#400 gamma=32'd4;row=32'd149;
#400 gamma=32'd5;row=32'd536;
#400 gamma=32'd5;row=32'd335;
#400 gamma=32'd5;row=32'd407;
#400 gamma=32'd3;row=32'd107;
#400 gamma=32'd3;row=32'd371;
#400 gamma=32'd3;row=32'd290;
#400 gamma=32'd1;row=32'd233;
#400 gamma=32'd5;row=32'd64;
#400 gamma=32'd2;row=32'd289;
#400 gamma=32'd2;row=32'd315;
#400 gamma=32'd5;row=32'd384;
#400 gamma=32'd4;row=32'd539;
#400 gamma=32'd1;row=32'd249;
#400 gamma=32'd1;row=32'd184;
#400 gamma=32'd5;row=32'd144;
#400 gamma=32'd1;row=32'd353;
#400 gamma=32'd3;row=32'd543;
#400 gamma=32'd5;row=32'd282;
#400 gamma=32'd4;row=32'd368;
#400 gamma=32'd4;row=32'd515;
#400 gamma=32'd5;row=32'd361;
#400 gamma=32'd2;row=32'd222;
#400 gamma=32'd3;row=32'd266;
#400 gamma=32'd3;row=32'd139;
#400 gamma=32'd5;row=32'd242;
#400 gamma=32'd5;row=32'd257;
#400 gamma=32'd4;row=32'd263;
#400 gamma=32'd1;row=32'd456;
#400 gamma=32'd1;row=32'd526;
#400 gamma=32'd2;row=32'd315;
#400 gamma=32'd4;row=32'd501;
#400 gamma=32'd1;row=32'd511;
#400 gamma=32'd2;row=32'd131;
#400 gamma=32'd4;row=32'd454;
#400 gamma=32'd4;row=32'd248;
#400 gamma=32'd2;row=32'd547;
#400 gamma=32'd2;row=32'd102;
#400 gamma=32'd1;row=32'd502;
#400 gamma=32'd4;row=32'd425;
#400 gamma=32'd2;row=32'd477;
#400 gamma=32'd1;row=32'd321;
#400 gamma=32'd4;row=32'd500;
#400 gamma=32'd2;row=32'd311;
#400 gamma=32'd3;row=32'd93;
#400 gamma=32'd5;row=32'd32;
#400 gamma=32'd3;row=32'd464;
#400 gamma=32'd5;row=32'd201;
#400 gamma=32'd2;row=32'd558;
#400 gamma=32'd4;row=32'd158;
#400 gamma=32'd4;row=32'd500;
#400 gamma=32'd4;row=32'd317;
#400 gamma=32'd2;row=32'd103;
#400 gamma=32'd3;row=32'd3;
#400 gamma=32'd2;row=32'd117;
#400 gamma=32'd2;row=32'd146;
#400 gamma=32'd4;row=32'd401;
#400 gamma=32'd4;row=32'd344;
#400 gamma=32'd3;row=32'd461;
#400 gamma=32'd5;row=32'd554;
#400 gamma=32'd2;row=32'd233;
#400 gamma=32'd1;row=32'd152;
#400 gamma=32'd2;row=32'd183;
#400 gamma=32'd2;row=32'd229;
#400 gamma=32'd4;row=32'd392;
#400 gamma=32'd4;row=32'd408;
#400 gamma=32'd4;row=32'd480;
#400 gamma=32'd4;row=32'd495;
#400 gamma=32'd2;row=32'd147;
#400 gamma=32'd1;row=32'd48;
#400 gamma=32'd1;row=32'd26;
#400 gamma=32'd3;row=32'd3;
#400 gamma=32'd4;row=32'd453;
#400 gamma=32'd5;row=32'd201;
#400 gamma=32'd5;row=32'd110;
#400 gamma=32'd2;row=32'd16;
#400 gamma=32'd5;row=32'd244;
#400 gamma=32'd3;row=32'd343;
#400 gamma=32'd4;row=32'd414;
#400 gamma=32'd5;row=32'd53;
#400 gamma=32'd3;row=32'd434;
#400 gamma=32'd1;row=32'd237;
#400 gamma=32'd3;row=32'd316;
#400 gamma=32'd2;row=32'd410;
#400 gamma=32'd1;row=32'd460;
#400 gamma=32'd1;row=32'd87;
#400 gamma=32'd5;row=32'd228;
#400 gamma=32'd3;row=32'd430;
#400 gamma=32'd5;row=32'd68;
#400 gamma=32'd4;row=32'd103;
#400 gamma=32'd1;row=32'd436;
#400 gamma=32'd4;row=32'd281;
#400 gamma=32'd3;row=32'd5;
#400 gamma=32'd2;row=32'd471;
#400 gamma=32'd1;row=32'd536;
#400 gamma=32'd5;row=32'd212;
#400 gamma=32'd4;row=32'd358;
#400 gamma=32'd4;row=32'd139;
#400 gamma=32'd5;row=32'd441;
#400 gamma=32'd2;row=32'd30;
#400 gamma=32'd1;row=32'd477;
#400 gamma=32'd1;row=32'd204;
#400 gamma=32'd2;row=32'd559;
#400 gamma=32'd5;row=32'd370;
#400 gamma=32'd2;row=32'd552;
#400 gamma=32'd5;row=32'd185;
#400 gamma=32'd2;row=32'd213;
#400 gamma=32'd5;row=32'd477;
#400 gamma=32'd5;row=32'd525;
#400 gamma=32'd1;row=32'd536;
#400 gamma=32'd1;row=32'd350;
#400 gamma=32'd1;row=32'd530;
#400 gamma=32'd4;row=32'd512;
#400 gamma=32'd2;row=32'd458;
#400 gamma=32'd3;row=32'd14;
#400 gamma=32'd1;row=32'd177;
#400 gamma=32'd1;row=32'd179;
#400 gamma=32'd3;row=32'd339;
#400 gamma=32'd2;row=32'd179;
#400 gamma=32'd3;row=32'd523;
#400 gamma=32'd4;row=32'd237;
#400 gamma=32'd5;row=32'd107;
#400 gamma=32'd1;row=32'd486;
#400 gamma=32'd1;row=32'd49;
#400 gamma=32'd5;row=32'd241;
#400 gamma=32'd3;row=32'd23;
#400 gamma=32'd5;row=32'd511;
#400 gamma=32'd3;row=32'd306;
#400 gamma=32'd3;row=32'd143;
#400 gamma=32'd1;row=32'd435;
#400 gamma=32'd2;row=32'd410;
#400 gamma=32'd2;row=32'd458;
#400 gamma=32'd4;row=32'd445;
#400 gamma=32'd3;row=32'd433;
#400 gamma=32'd2;row=32'd208;
#400 gamma=32'd5;row=32'd124;
#400 gamma=32'd1;row=32'd47;
#400 gamma=32'd5;row=32'd127;
#400 gamma=32'd1;row=32'd118;
#400 gamma=32'd3;row=32'd18;
#400 gamma=32'd2;row=32'd213;
#400 gamma=32'd1;row=32'd460;
#400 gamma=32'd4;row=32'd521;
#400 gamma=32'd3;row=32'd299;
#400 gamma=32'd5;row=32'd95;
#400 gamma=32'd2;row=32'd204;
#400 gamma=32'd3;row=32'd549;
#400 gamma=32'd4;row=32'd544;
#400 gamma=32'd1;row=32'd217;
#400 gamma=32'd4;row=32'd422;
#400 gamma=32'd5;row=32'd139;
#400 gamma=32'd3;row=32'd543;
#400 gamma=32'd2;row=32'd474;
#400 gamma=32'd3;row=32'd103;
#400 gamma=32'd3;row=32'd514;
#400 gamma=32'd1;row=32'd22;
#400 gamma=32'd5;row=32'd556;
#400 gamma=32'd1;row=32'd99;
#400 gamma=32'd4;row=32'd414;
#400 gamma=32'd2;row=32'd552;
#400 gamma=32'd1;row=32'd271;
#400 gamma=32'd3;row=32'd237;
#400 gamma=32'd1;row=32'd235;
#400 gamma=32'd1;row=32'd352;
#400 gamma=32'd5;row=32'd51;
#400 gamma=32'd3;row=32'd62;
#400 gamma=32'd4;row=32'd1;
#400 gamma=32'd1;row=32'd325;
#400 gamma=32'd1;row=32'd341;
#400 gamma=32'd1;row=32'd86;
#400 gamma=32'd2;row=32'd37;
#400 gamma=32'd4;row=32'd363;
#400 gamma=32'd4;row=32'd57;
#400 gamma=32'd3;row=32'd402;
#400 gamma=32'd2;row=32'd48;
#400 gamma=32'd1;row=32'd138;
#400 gamma=32'd2;row=32'd479;
#400 gamma=32'd3;row=32'd394;
#400 gamma=32'd5;row=32'd272;
#400 gamma=32'd5;row=32'd193;
#400 gamma=32'd1;row=32'd247;
#400 gamma=32'd1;row=32'd477;
#400 gamma=32'd4;row=32'd343;
#400 gamma=32'd2;row=32'd157;
#400 gamma=32'd4;row=32'd129;
#400 gamma=32'd5;row=32'd98;
#400 gamma=32'd2;row=32'd355;
#400 gamma=32'd5;row=32'd544;
#400 gamma=32'd4;row=32'd494;
#400 gamma=32'd2;row=32'd497;
#400 gamma=32'd5;row=32'd539;
#400 gamma=32'd1;row=32'd55;
#400 gamma=32'd2;row=32'd229;
#400 gamma=32'd5;row=32'd154;
#400 gamma=32'd2;row=32'd62;
#400 gamma=32'd3;row=32'd429;
#400 gamma=32'd2;row=32'd385;
#400 gamma=32'd3;row=32'd49;
#400 gamma=32'd4;row=32'd122;
#400 gamma=32'd1;row=32'd171;
#400 gamma=32'd4;row=32'd320;
#400 gamma=32'd1;row=32'd46;
#400 gamma=32'd4;row=32'd237;
#400 gamma=32'd4;row=32'd210;
#400 gamma=32'd5;row=32'd457;
#400 gamma=32'd1;row=32'd475;
#400 gamma=32'd3;row=32'd54;
#400 gamma=32'd5;row=32'd47;
#400 gamma=32'd4;row=32'd496;
#400 gamma=32'd1;row=32'd310;
#400 gamma=32'd1;row=32'd204;
#400 gamma=32'd1;row=32'd62;
#400 gamma=32'd1;row=32'd511;
#400 gamma=32'd1;row=32'd118;
#400 gamma=32'd3;row=32'd551;
#400 gamma=32'd4;row=32'd297;
#400 gamma=32'd5;row=32'd76;
#400 gamma=32'd2;row=32'd277;
#400 gamma=32'd3;row=32'd130;
#400 gamma=32'd1;row=32'd233;
#400 gamma=32'd1;row=32'd138;
#400 gamma=32'd1;row=32'd428;
#400 gamma=32'd5;row=32'd90;
#400 gamma=32'd3;row=32'd387;
#400 gamma=32'd1;row=32'd400;
#400 gamma=32'd4;row=32'd51;
#400 gamma=32'd2;row=32'd34;
#400 gamma=32'd3;row=32'd51;
#400 gamma=32'd1;row=32'd184;
#400 gamma=32'd4;row=32'd417;
#400 gamma=32'd1;row=32'd242;
#400 gamma=32'd2;row=32'd8;
#400 gamma=32'd4;row=32'd203;
#400 gamma=32'd4;row=32'd384;
#400 gamma=32'd1;row=32'd172;
#400 gamma=32'd5;row=32'd363;
#400 gamma=32'd2;row=32'd227;
#400 gamma=32'd1;row=32'd297;
#400 gamma=32'd5;row=32'd176;
#400 gamma=32'd5;row=32'd381;
#400 gamma=32'd3;row=32'd39;
#400 gamma=32'd5;row=32'd506;
#400 gamma=32'd4;row=32'd295;
#400 gamma=32'd3;row=32'd6;
#400 gamma=32'd1;row=32'd214;
#400 gamma=32'd2;row=32'd308;
#400 gamma=32'd5;row=32'd269;
#400 gamma=32'd5;row=32'd327;
#400 gamma=32'd5;row=32'd332;
#400 gamma=32'd2;row=32'd139;
#400 gamma=32'd4;row=32'd434;
#400 gamma=32'd4;row=32'd281;
#400 gamma=32'd3;row=32'd493;
#400 gamma=32'd2;row=32'd508;
#400 gamma=32'd5;row=32'd300;
#400 gamma=32'd5;row=32'd10;
#400 gamma=32'd3;row=32'd214;
#400 gamma=32'd3;row=32'd221;
#400 gamma=32'd2;row=32'd23;
#400 gamma=32'd3;row=32'd428;
#400 gamma=32'd4;row=32'd517;
#400 gamma=32'd3;row=32'd289;
#400 gamma=32'd5;row=32'd534;
#400 gamma=32'd3;row=32'd300;
#400 gamma=32'd2;row=32'd512;
#400 gamma=32'd5;row=32'd40;
#400 gamma=32'd4;row=32'd241;
#400 gamma=32'd4;row=32'd515;
#400 gamma=32'd4;row=32'd118;
#400 gamma=32'd1;row=32'd320;
#400 gamma=32'd2;row=32'd279;
#400 gamma=32'd4;row=32'd486;
#400 gamma=32'd4;row=32'd210;
#400 gamma=32'd3;row=32'd221;
#400 gamma=32'd4;row=32'd431;
#400 gamma=32'd1;row=32'd167;
#400 gamma=32'd1;row=32'd42;
#400 gamma=32'd4;row=32'd444;
#400 gamma=32'd2;row=32'd204;
#400 gamma=32'd3;row=32'd181;
#400 gamma=32'd4;row=32'd183;
#400 gamma=32'd5;row=32'd273;
#400 gamma=32'd3;row=32'd308;
#400 gamma=32'd5;row=32'd356;
#400 gamma=32'd1;row=32'd532;
#400 gamma=32'd4;row=32'd465;
#400 gamma=32'd2;row=32'd290;
#400 gamma=32'd4;row=32'd422;
#400 gamma=32'd1;row=32'd305;
#400 gamma=32'd1;row=32'd507;
#400 gamma=32'd5;row=32'd489;
#400 gamma=32'd4;row=32'd284;
#400 gamma=32'd3;row=32'd306;
#400 gamma=32'd5;row=32'd97;
#400 gamma=32'd3;row=32'd428;
#400 gamma=32'd1;row=32'd448;
#400 gamma=32'd5;row=32'd3;
#400 gamma=32'd2;row=32'd559;
#400 gamma=32'd2;row=32'd110;
#400 gamma=32'd1;row=32'd414;
#400 gamma=32'd3;row=32'd246;
#400 gamma=32'd3;row=32'd135;
#400 gamma=32'd5;row=32'd137;
#400 gamma=32'd4;row=32'd424;
#400 gamma=32'd5;row=32'd495;
#400 gamma=32'd1;row=32'd558;
#400 gamma=32'd4;row=32'd268;
#400 gamma=32'd3;row=32'd408;
#400 gamma=32'd1;row=32'd443;
#400 gamma=32'd5;row=32'd204;
#400 gamma=32'd2;row=32'd458;
#400 gamma=32'd4;row=32'd113;
#400 gamma=32'd4;row=32'd470;
#400 gamma=32'd4;row=32'd442;
#400 gamma=32'd4;row=32'd115;
#400 gamma=32'd1;row=32'd281;
#400 gamma=32'd2;row=32'd540;
#400 gamma=32'd4;row=32'd28;
#400 gamma=32'd2;row=32'd346;
#400 gamma=32'd2;row=32'd62;
#400 gamma=32'd1;row=32'd479;
#400 gamma=32'd1;row=32'd531;
#400 gamma=32'd2;row=32'd478;
#400 gamma=32'd1;row=32'd151;
#400 gamma=32'd5;row=32'd486;
#400 gamma=32'd1;row=32'd184;
#400 gamma=32'd4;row=32'd268;
#400 gamma=32'd1;row=32'd296;
#400 gamma=32'd5;row=32'd8;
#400 gamma=32'd5;row=32'd476;
#400 gamma=32'd4;row=32'd182;
#400 gamma=32'd4;row=32'd439;
#400 gamma=32'd5;row=32'd183;
#400 gamma=32'd5;row=32'd513;
#400 gamma=32'd1;row=32'd534;
#400 gamma=32'd4;row=32'd231;
#400 gamma=32'd2;row=32'd127;
#400 gamma=32'd3;row=32'd373;
#400 gamma=32'd3;row=32'd160;
#400 gamma=32'd4;row=32'd142;
#400 gamma=32'd4;row=32'd437;
#400 gamma=32'd4;row=32'd0;
#400 gamma=32'd3;row=32'd442;
#400 gamma=32'd3;row=32'd448;
#400 gamma=32'd1;row=32'd405;
#400 gamma=32'd4;row=32'd31;
#400 gamma=32'd4;row=32'd367;
#400 gamma=32'd1;row=32'd511;
#400 gamma=32'd2;row=32'd239;
#400 gamma=32'd2;row=32'd238;
#400 gamma=32'd1;row=32'd457;
#400 gamma=32'd4;row=32'd218;
#400 gamma=32'd3;row=32'd187;
#400 gamma=32'd2;row=32'd500;
#400 gamma=32'd2;row=32'd39;
#400 gamma=32'd2;row=32'd526;
#400 gamma=32'd2;row=32'd297;
#400 gamma=32'd5;row=32'd195;
#400 gamma=32'd5;row=32'd285;
#400 gamma=32'd5;row=32'd552;
#400 gamma=32'd4;row=32'd195;
#400 gamma=32'd5;row=32'd58;
#400 gamma=32'd2;row=32'd178;
#400 gamma=32'd5;row=32'd20;
#400 gamma=32'd2;row=32'd412;
#400 gamma=32'd4;row=32'd487;
#400 gamma=32'd1;row=32'd305;
#400 gamma=32'd1;row=32'd51;
#400 gamma=32'd5;row=32'd348;
#400 gamma=32'd4;row=32'd265;
#400 gamma=32'd3;row=32'd492;
#400 gamma=32'd4;row=32'd197;
#400 gamma=32'd3;row=32'd31;
#400 gamma=32'd4;row=32'd541;
#400 gamma=32'd5;row=32'd221;
#400 gamma=32'd1;row=32'd54;
#400 gamma=32'd3;row=32'd32;
#400 gamma=32'd2;row=32'd558;
#400 gamma=32'd2;row=32'd399;
#400 gamma=32'd5;row=32'd60;
#400 gamma=32'd5;row=32'd103;
#400 gamma=32'd2;row=32'd433;
#400 gamma=32'd2;row=32'd19;
#400 gamma=32'd4;row=32'd82;
#400 gamma=32'd5;row=32'd526;
#400 gamma=32'd5;row=32'd120;
#400 gamma=32'd5;row=32'd12;
#400 gamma=32'd2;row=32'd146;
#400 gamma=32'd5;row=32'd434;
#400 gamma=32'd5;row=32'd382;
#400 gamma=32'd4;row=32'd74;
#400 gamma=32'd4;row=32'd529;
#400 gamma=32'd3;row=32'd67;
#400 gamma=32'd1;row=32'd39;
#400 gamma=32'd5;row=32'd270;
#400 gamma=32'd5;row=32'd364;
#400 gamma=32'd3;row=32'd124;
#400 gamma=32'd3;row=32'd138;
#400 gamma=32'd2;row=32'd434;
#400 gamma=32'd3;row=32'd79;
#400 gamma=32'd1;row=32'd348;
#400 gamma=32'd5;row=32'd142;
#400 gamma=32'd2;row=32'd456;
#400 gamma=32'd5;row=32'd8;
#400 gamma=32'd5;row=32'd260;
#400 gamma=32'd5;row=32'd38;
#400 gamma=32'd5;row=32'd240;
#400 gamma=32'd2;row=32'd128;
#400 gamma=32'd2;row=32'd395;
#400 gamma=32'd3;row=32'd290;
#400 gamma=32'd1;row=32'd37;
#400 gamma=32'd1;row=32'd226;
#400 gamma=32'd5;row=32'd216;
#400 gamma=32'd1;row=32'd213;
#400 gamma=32'd1;row=32'd397;
#400 gamma=32'd4;row=32'd280;
#400 gamma=32'd1;row=32'd182;
#400 gamma=32'd5;row=32'd519;
#400 gamma=32'd5;row=32'd164;
#400 gamma=32'd1;row=32'd454;
#400 gamma=32'd2;row=32'd227;
#400 gamma=32'd3;row=32'd365;
#400 gamma=32'd5;row=32'd473;
#400 gamma=32'd3;row=32'd501;
#400 gamma=32'd4;row=32'd401;
#400 gamma=32'd5;row=32'd317;
#400 gamma=32'd3;row=32'd464;
#400 gamma=32'd2;row=32'd467;
#400 gamma=32'd2;row=32'd192;
#400 gamma=32'd3;row=32'd355;
#400 gamma=32'd2;row=32'd504;
#400 gamma=32'd4;row=32'd100;
#400 gamma=32'd4;row=32'd375;
#400 gamma=32'd5;row=32'd499;
#400 gamma=32'd1;row=32'd214;
#400 gamma=32'd3;row=32'd305;
#400 gamma=32'd5;row=32'd69;
#400 gamma=32'd3;row=32'd99;
#400 gamma=32'd3;row=32'd111;
#400 gamma=32'd5;row=32'd236;
#400 gamma=32'd2;row=32'd350;
#400 gamma=32'd1;row=32'd506;
#400 gamma=32'd5;row=32'd367;
#400 gamma=32'd4;row=32'd88;
#400 gamma=32'd4;row=32'd181;
#400 gamma=32'd1;row=32'd81;
#400 gamma=32'd3;row=32'd507;
#400 gamma=32'd5;row=32'd279;
#400 gamma=32'd3;row=32'd510;
#400 gamma=32'd2;row=32'd387;
#400 gamma=32'd4;row=32'd524;
#400 gamma=32'd4;row=32'd227;
#400 gamma=32'd2;row=32'd291;
#400 gamma=32'd5;row=32'd229;
#400 gamma=32'd5;row=32'd398;
#400 gamma=32'd3;row=32'd343;
#400 gamma=32'd2;row=32'd321;
#400 gamma=32'd4;row=32'd508;
#400 gamma=32'd3;row=32'd217;
#400 gamma=32'd3;row=32'd469;
#400 gamma=32'd1;row=32'd375;
#400 gamma=32'd2;row=32'd229;
#400 gamma=32'd5;row=32'd306;
#400 gamma=32'd1;row=32'd308;
#400 gamma=32'd3;row=32'd441;
#400 gamma=32'd4;row=32'd232;
#400 gamma=32'd2;row=32'd291;
#400 gamma=32'd1;row=32'd85;
#400 gamma=32'd2;row=32'd524;
#400 gamma=32'd5;row=32'd297;
#400 gamma=32'd1;row=32'd45;
#400 gamma=32'd1;row=32'd409;
#400 gamma=32'd4;row=32'd394;
#400 gamma=32'd4;row=32'd162;
#400 gamma=32'd5;row=32'd396;
#400 gamma=32'd5;row=32'd255;
#400 gamma=32'd4;row=32'd182;
#400 gamma=32'd5;row=32'd157;
#400 gamma=32'd4;row=32'd9;
#400 gamma=32'd3;row=32'd407;
#400 gamma=32'd5;row=32'd120;
#400 gamma=32'd2;row=32'd420;
#400 gamma=32'd4;row=32'd415;
#400 gamma=32'd1;row=32'd314;
#400 gamma=32'd5;row=32'd36;
#400 gamma=32'd5;row=32'd167;
#400 gamma=32'd4;row=32'd224;
#400 gamma=32'd1;row=32'd505;
#400 gamma=32'd5;row=32'd340;
#400 gamma=32'd2;row=32'd303;
#400 gamma=32'd4;row=32'd341;
#400 gamma=32'd3;row=32'd348;
#400 gamma=32'd5;row=32'd162;
#400 gamma=32'd5;row=32'd480;
#400 gamma=32'd3;row=32'd302;
#400 gamma=32'd3;row=32'd304;
#400 gamma=32'd3;row=32'd79;
#400 gamma=32'd2;row=32'd89;
#400 gamma=32'd1;row=32'd470;
#400 gamma=32'd2;row=32'd489;
#400 gamma=32'd4;row=32'd223;
#400 gamma=32'd1;row=32'd95;
#400 gamma=32'd2;row=32'd510;
#400 gamma=32'd5;row=32'd454;
#400 gamma=32'd3;row=32'd200;
#400 gamma=32'd4;row=32'd308;
#400 gamma=32'd4;row=32'd280;
#400 gamma=32'd2;row=32'd6;
#400 gamma=32'd5;row=32'd28;
#400 gamma=32'd5;row=32'd18;
#400 gamma=32'd4;row=32'd348;
#400 gamma=32'd5;row=32'd526;
#400 gamma=32'd3;row=32'd261;
#400 gamma=32'd4;row=32'd315;
#400 gamma=32'd4;row=32'd479;
#400 gamma=32'd3;row=32'd380;
#400 gamma=32'd3;row=32'd287;
#400 gamma=32'd1;row=32'd399;
#400 gamma=32'd4;row=32'd248;
#400 gamma=32'd4;row=32'd227;
#400 gamma=32'd4;row=32'd89;
#400 gamma=32'd1;row=32'd212;
#400 gamma=32'd1;row=32'd497;
#400 gamma=32'd1;row=32'd329;
#400 gamma=32'd3;row=32'd139;
#400 gamma=32'd5;row=32'd213;
#400 gamma=32'd3;row=32'd307;
#400 gamma=32'd2;row=32'd180;
#400 gamma=32'd2;row=32'd397;
#400 gamma=32'd1;row=32'd441;
#400 gamma=32'd5;row=32'd387;
#400 gamma=32'd3;row=32'd391;
#400 gamma=32'd5;row=32'd184;
#400 gamma=32'd3;row=32'd336;
#400 gamma=32'd1;row=32'd254;
#400 gamma=32'd1;row=32'd550;
#400 gamma=32'd5;row=32'd57;
#400 gamma=32'd1;row=32'd188;
#400 gamma=32'd4;row=32'd286;
#400 gamma=32'd5;row=32'd175;
#400 gamma=32'd3;row=32'd517;
#400 gamma=32'd3;row=32'd447;
#400 gamma=32'd2;row=32'd164;
#400 gamma=32'd1;row=32'd335;
#400 gamma=32'd5;row=32'd208;
#400 gamma=32'd3;row=32'd306;
#400 gamma=32'd5;row=32'd121;
#400 gamma=32'd4;row=32'd493;
#400 gamma=32'd2;row=32'd304;
#400 gamma=32'd1;row=32'd1;
#400 gamma=32'd4;row=32'd307;
#400 gamma=32'd2;row=32'd189;
#400 gamma=32'd1;row=32'd559;
#400 gamma=32'd2;row=32'd325;
#400 gamma=32'd1;row=32'd248;
#400 gamma=32'd3;row=32'd205;
#400 gamma=32'd4;row=32'd157;
#400 gamma=32'd2;row=32'd541;
#400 gamma=32'd3;row=32'd143;
#400 gamma=32'd5;row=32'd173;
#400 gamma=32'd2;row=32'd141;
#400 gamma=32'd4;row=32'd212;
#400 gamma=32'd3;row=32'd555;
#400 gamma=32'd3;row=32'd401;
#400 gamma=32'd1;row=32'd371;
#400 gamma=32'd4;row=32'd264;
#400 gamma=32'd3;row=32'd354;
#400 gamma=32'd1;row=32'd539;
#400 gamma=32'd4;row=32'd468;
#400 gamma=32'd4;row=32'd226;
#400 gamma=32'd4;row=32'd493;
#400 gamma=32'd4;row=32'd240;
#400 gamma=32'd1;row=32'd287;
#400 gamma=32'd5;row=32'd20;
#400 gamma=32'd1;row=32'd256;
#400 gamma=32'd5;row=32'd295;
#400 gamma=32'd1;row=32'd403;
#400 gamma=32'd2;row=32'd478;
#400 gamma=32'd2;row=32'd475;
#400 gamma=32'd2;row=32'd524;
#400 gamma=32'd1;row=32'd186;
#400 gamma=32'd4;row=32'd231;
#400 gamma=32'd1;row=32'd504;
#400 gamma=32'd5;row=32'd533;
#400 gamma=32'd3;row=32'd342;
#400 gamma=32'd1;row=32'd450;
#400 gamma=32'd2;row=32'd139;
#400 gamma=32'd1;row=32'd224;
#400 gamma=32'd2;row=32'd16;
#400 gamma=32'd2;row=32'd165;
#400 gamma=32'd1;row=32'd272;
#400 gamma=32'd5;row=32'd33;
#400 gamma=32'd2;row=32'd35;
#400 gamma=32'd5;row=32'd17;
#400 gamma=32'd2;row=32'd16;
#400 gamma=32'd5;row=32'd557;
#400 gamma=32'd3;row=32'd17;
#400 gamma=32'd1;row=32'd207;
#400 gamma=32'd3;row=32'd250;
#400 gamma=32'd2;row=32'd427;
#400 gamma=32'd4;row=32'd405;
#400 gamma=32'd1;row=32'd475;
#400 gamma=32'd4;row=32'd465;
#400 gamma=32'd1;row=32'd475;
#400 gamma=32'd3;row=32'd503;
#400 gamma=32'd5;row=32'd451;
#400 gamma=32'd4;row=32'd517;
#400 gamma=32'd3;row=32'd0;
#400 gamma=32'd5;row=32'd415;
#400 gamma=32'd4;row=32'd195;
#400 gamma=32'd1;row=32'd252;
#400 gamma=32'd5;row=32'd11;
#400 gamma=32'd4;row=32'd236;
#400 gamma=32'd2;row=32'd436;
#400 gamma=32'd2;row=32'd414;
#400 gamma=32'd1;row=32'd526;
#400 gamma=32'd2;row=32'd427;
#400 gamma=32'd1;row=32'd511;
#400 gamma=32'd3;row=32'd146;
#400 gamma=32'd2;row=32'd185;
#400 gamma=32'd3;row=32'd60;
#400 gamma=32'd2;row=32'd321;
#400 gamma=32'd3;row=32'd275;
#400 gamma=32'd5;row=32'd443;
#400 gamma=32'd2;row=32'd371;
#400 gamma=32'd2;row=32'd37;
#400 gamma=32'd3;row=32'd406;
#400 gamma=32'd5;row=32'd555;
#400 gamma=32'd4;row=32'd172;
#400 gamma=32'd1;row=32'd276;
#400 gamma=32'd5;row=32'd167;
#400 gamma=32'd2;row=32'd315;
#400 gamma=32'd4;row=32'd184;
#400 gamma=32'd5;row=32'd84;
#400 gamma=32'd5;row=32'd369;
#400 gamma=32'd4;row=32'd539;
#400 gamma=32'd3;row=32'd536;
#400 gamma=32'd3;row=32'd56;
#400 gamma=32'd2;row=32'd394;
#400 gamma=32'd4;row=32'd56;
#400 gamma=32'd5;row=32'd125;
#400 gamma=32'd4;row=32'd438;
#400 gamma=32'd1;row=32'd149;
#400 gamma=32'd3;row=32'd546;
#400 gamma=32'd3;row=32'd100;
#400 gamma=32'd5;row=32'd521;
#400 gamma=32'd3;row=32'd29;
#400 gamma=32'd1;row=32'd347;
#400 gamma=32'd1;row=32'd86;
#400 gamma=32'd5;row=32'd537;
#400 gamma=32'd1;row=32'd411;
#400 gamma=32'd1;row=32'd477;
#400 gamma=32'd3;row=32'd533;
#400 gamma=32'd4;row=32'd518;
#400 gamma=32'd5;row=32'd434;
#400 gamma=32'd3;row=32'd38;
#400 gamma=32'd1;row=32'd50;
#400 gamma=32'd3;row=32'd364;
#400 gamma=32'd1;row=32'd193;
#400 gamma=32'd1;row=32'd110;
#400 gamma=32'd2;row=32'd243;
#400 gamma=32'd3;row=32'd380;
#400 gamma=32'd5;row=32'd95;
#400 gamma=32'd5;row=32'd20;
#400 gamma=32'd2;row=32'd144;
#400 gamma=32'd4;row=32'd404;
#400 gamma=32'd3;row=32'd460;
#400 gamma=32'd5;row=32'd448;
#400 gamma=32'd3;row=32'd79;
#400 gamma=32'd1;row=32'd74;
#400 gamma=32'd4;row=32'd285;
#400 gamma=32'd2;row=32'd558;
#400 gamma=32'd5;row=32'd523;
#400 gamma=32'd5;row=32'd382;
#400 gamma=32'd2;row=32'd63;
#400 gamma=32'd1;row=32'd289;
#400 gamma=32'd5;row=32'd45;
#400 gamma=32'd2;row=32'd362;
#400 gamma=32'd2;row=32'd73;
#400 gamma=32'd2;row=32'd206;
#400 gamma=32'd2;row=32'd348;
#400 gamma=32'd2;row=32'd327;
#400 gamma=32'd3;row=32'd536;
#400 gamma=32'd2;row=32'd175;
#400 gamma=32'd4;row=32'd309;
#400 gamma=32'd2;row=32'd390;
#400 gamma=32'd2;row=32'd109;
#400 gamma=32'd1;row=32'd203;
#400 gamma=32'd3;row=32'd236;
#400 gamma=32'd2;row=32'd93;
#400 gamma=32'd5;row=32'd130;
#400 gamma=32'd4;row=32'd297;
#400 gamma=32'd3;row=32'd320;
#400 gamma=32'd2;row=32'd472;
#400 gamma=32'd1;row=32'd468;
#400 gamma=32'd5;row=32'd294;
#400 gamma=32'd5;row=32'd131;
#400 gamma=32'd3;row=32'd532;
#400 gamma=32'd5;row=32'd219;
#400 gamma=32'd5;row=32'd376;
#400 gamma=32'd1;row=32'd111;
#400 gamma=32'd4;row=32'd80;
#400 gamma=32'd1;row=32'd313;
#400 gamma=32'd2;row=32'd519;
#400 gamma=32'd5;row=32'd237;
#400 gamma=32'd1;row=32'd67;
#400 gamma=32'd5;row=32'd448;
#400 gamma=32'd1;row=32'd222;
#400 gamma=32'd4;row=32'd416;
#400 gamma=32'd1;row=32'd144;
#400 gamma=32'd1;row=32'd17;
#400 gamma=32'd2;row=32'd87;
#400 gamma=32'd5;row=32'd96;
#400 gamma=32'd2;row=32'd248;
#400 gamma=32'd2;row=32'd288;
#400 gamma=32'd4;row=32'd443;
#400 gamma=32'd1;row=32'd47;
#400 gamma=32'd3;row=32'd324;
#400 gamma=32'd2;row=32'd398;
#400 gamma=32'd3;row=32'd306;
#400 gamma=32'd5;row=32'd9;
#400 gamma=32'd3;row=32'd29;
#400 gamma=32'd3;row=32'd339;
#400 gamma=32'd4;row=32'd403;
#400 gamma=32'd4;row=32'd205;
#400 gamma=32'd3;row=32'd208;
#400 gamma=32'd1;row=32'd138;
#400 gamma=32'd5;row=32'd519;
#400 gamma=32'd5;row=32'd11;
#400 gamma=32'd2;row=32'd216;
#400 gamma=32'd4;row=32'd72;
#400 gamma=32'd1;row=32'd358;
#400 gamma=32'd1;row=32'd462;
#400 gamma=32'd5;row=32'd383;
#400 gamma=32'd5;row=32'd209;
#400 gamma=32'd1;row=32'd286;
#400 gamma=32'd4;row=32'd74;
#400 gamma=32'd3;row=32'd349;
#400 gamma=32'd4;row=32'd389;
#400 gamma=32'd5;row=32'd422;
#400 gamma=32'd4;row=32'd119;
#400 gamma=32'd1;row=32'd357;
#400 gamma=32'd3;row=32'd241;
#400 gamma=32'd1;row=32'd486;
#400 gamma=32'd3;row=32'd10;
#400 gamma=32'd2;row=32'd474;
#400 gamma=32'd5;row=32'd152;
#400 gamma=32'd3;row=32'd375;
#400 gamma=32'd1;row=32'd116;
#400 gamma=32'd5;row=32'd223;
#400 gamma=32'd4;row=32'd127;
#400 gamma=32'd5;row=32'd486;
#400 gamma=32'd3;row=32'd529;
#400 gamma=32'd2;row=32'd119;
#400 gamma=32'd1;row=32'd366;
#400 gamma=32'd1;row=32'd207;
#400 gamma=32'd4;row=32'd349;
#400 gamma=32'd3;row=32'd93;
#400 gamma=32'd5;row=32'd168;
#400 gamma=32'd3;row=32'd35;
#400 gamma=32'd2;row=32'd541;
#400 gamma=32'd1;row=32'd340;
#400 gamma=32'd4;row=32'd273;
#400 gamma=32'd4;row=32'd92;
#400 gamma=32'd1;row=32'd47;
#400 gamma=32'd4;row=32'd254;
#400 gamma=32'd4;row=32'd59;
#400 gamma=32'd5;row=32'd445;
#400 gamma=32'd1;row=32'd334;
#400 gamma=32'd2;row=32'd9;
#400 gamma=32'd4;row=32'd128;
#400 gamma=32'd1;row=32'd432;
#400 gamma=32'd4;row=32'd129;
#400 gamma=32'd3;row=32'd126;
#400 gamma=32'd1;row=32'd48;
#400 gamma=32'd5;row=32'd144;
#400 gamma=32'd1;row=32'd248;
#400 gamma=32'd1;row=32'd465;
#400 gamma=32'd4;row=32'd110;
#400 gamma=32'd2;row=32'd97;
#400 gamma=32'd1;row=32'd337;
#400 gamma=32'd4;row=32'd400;
#400 gamma=32'd1;row=32'd406;
#400 gamma=32'd5;row=32'd354;
#400 gamma=32'd5;row=32'd286;
#400 gamma=32'd2;row=32'd176;
#400 gamma=32'd1;row=32'd312;
#400 gamma=32'd4;row=32'd368;
#400 gamma=32'd5;row=32'd250;
#400 gamma=32'd5;row=32'd90;
#400 gamma=32'd4;row=32'd79;
#400 gamma=32'd2;row=32'd113;
#400 gamma=32'd4;row=32'd55;
#400 gamma=32'd4;row=32'd501;
#400 gamma=32'd3;row=32'd66;
#400 gamma=32'd3;row=32'd363;
#400 gamma=32'd5;row=32'd302;
#400 gamma=32'd1;row=32'd198;
#400 gamma=32'd3;row=32'd383;
#400 gamma=32'd3;row=32'd278;
#400 gamma=32'd4;row=32'd415;
#400 gamma=32'd3;row=32'd291;
#400 gamma=32'd2;row=32'd99;
#400 gamma=32'd4;row=32'd322;
#400 gamma=32'd5;row=32'd387;
#400 gamma=32'd1;row=32'd201;
#400 gamma=32'd1;row=32'd392;
#400 gamma=32'd4;row=32'd510;
#400 gamma=32'd3;row=32'd15;
#400 gamma=32'd2;row=32'd90;
#400 gamma=32'd2;row=32'd111;
#400 gamma=32'd4;row=32'd258;
#400 gamma=32'd3;row=32'd538;
#400 gamma=32'd1;row=32'd39;
#400 gamma=32'd5;row=32'd111;
#400 gamma=32'd4;row=32'd452;
#400 gamma=32'd5;row=32'd504;
#400 gamma=32'd4;row=32'd555;
#400 gamma=32'd5;row=32'd8;
#400 gamma=32'd2;row=32'd366;
#400 gamma=32'd5;row=32'd250;
#400 gamma=32'd4;row=32'd39;
#400 gamma=32'd5;row=32'd346;
#400 gamma=32'd2;row=32'd489;
#400 gamma=32'd1;row=32'd379;
#400 gamma=32'd1;row=32'd305;
#400 gamma=32'd2;row=32'd36;
#400 gamma=32'd1;row=32'd352;
#400 gamma=32'd1;row=32'd193;
#400 gamma=32'd3;row=32'd368;
#400 gamma=32'd3;row=32'd268;
#400 gamma=32'd5;row=32'd195;
#400 gamma=32'd1;row=32'd11;
#400 gamma=32'd5;row=32'd517;
#400 gamma=32'd2;row=32'd75;
#400 gamma=32'd4;row=32'd243;
#400 gamma=32'd1;row=32'd395;
#400 gamma=32'd1;row=32'd557;
#400 gamma=32'd4;row=32'd323;
#400 gamma=32'd5;row=32'd146;
#400 gamma=32'd1;row=32'd15;
#400 gamma=32'd2;row=32'd532;
#400 gamma=32'd5;row=32'd384;
#400 gamma=32'd4;row=32'd387;
#400 gamma=32'd1;row=32'd165;
#400 gamma=32'd2;row=32'd32;
#400 gamma=32'd2;row=32'd516;
#400 gamma=32'd5;row=32'd88;
#400 gamma=32'd5;row=32'd244;
#400 gamma=32'd4;row=32'd171;
#400 gamma=32'd4;row=32'd253;
#400 gamma=32'd3;row=32'd167;
#400 gamma=32'd5;row=32'd513;
#400 gamma=32'd3;row=32'd245;
#400 gamma=32'd1;row=32'd367;
#400 gamma=32'd5;row=32'd193;
#400 gamma=32'd4;row=32'd12;
#400 gamma=32'd1;row=32'd228;
#400 gamma=32'd5;row=32'd206;
#400 gamma=32'd2;row=32'd159;
#400 gamma=32'd4;row=32'd557;
#400 gamma=32'd5;row=32'd474;
#400 gamma=32'd3;row=32'd135;
#400 gamma=32'd1;row=32'd395;
#400 gamma=32'd5;row=32'd198;
#400 gamma=32'd4;row=32'd549;
#400 gamma=32'd2;row=32'd123;
#400 gamma=32'd4;row=32'd372;
#400 gamma=32'd4;row=32'd441;
#400 gamma=32'd5;row=32'd223;
#400 gamma=32'd3;row=32'd71;
#400 gamma=32'd2;row=32'd221;
#400 gamma=32'd3;row=32'd27;
#400 gamma=32'd1;row=32'd298;
#400 gamma=32'd3;row=32'd340;
#400 gamma=32'd1;row=32'd355;
#400 gamma=32'd5;row=32'd133;
#400 gamma=32'd3;row=32'd4;
#400 gamma=32'd5;row=32'd87;
#400 gamma=32'd1;row=32'd478;
#400 gamma=32'd5;row=32'd327;
#400 gamma=32'd5;row=32'd118;
#400 gamma=32'd2;row=32'd406;
#400 gamma=32'd2;row=32'd282;
#400 gamma=32'd2;row=32'd220;
#400 gamma=32'd5;row=32'd152;
#400 gamma=32'd4;row=32'd514;
#400 gamma=32'd2;row=32'd349;
#400 gamma=32'd2;row=32'd425;
#400 gamma=32'd2;row=32'd241;
#400 gamma=32'd4;row=32'd61;
#400 gamma=32'd2;row=32'd150;
#400 gamma=32'd5;row=32'd134;
#400 gamma=32'd5;row=32'd445;
#400 gamma=32'd2;row=32'd406;
#400 gamma=32'd2;row=32'd243;
#400 gamma=32'd2;row=32'd556;
#400 gamma=32'd1;row=32'd266;
#400 gamma=32'd3;row=32'd121;
#400 gamma=32'd5;row=32'd326;
#400 gamma=32'd4;row=32'd1;
#400 gamma=32'd2;row=32'd21;
#400 gamma=32'd4;row=32'd214;
#400 gamma=32'd4;row=32'd216;
#400 gamma=32'd4;row=32'd411;
#400 gamma=32'd3;row=32'd410;
#400 gamma=32'd1;row=32'd192;
#400 gamma=32'd3;row=32'd264;
#400 gamma=32'd2;row=32'd201;
#400 gamma=32'd2;row=32'd545;
#400 gamma=32'd1;row=32'd13;
#400 gamma=32'd1;row=32'd487;
#400 gamma=32'd2;row=32'd167;
#400 gamma=32'd4;row=32'd9;
#400 gamma=32'd2;row=32'd15;
#400 gamma=32'd4;row=32'd399;
#400 gamma=32'd1;row=32'd381;
#400 gamma=32'd3;row=32'd64;
#400 gamma=32'd5;row=32'd485;
#400 gamma=32'd4;row=32'd308;
#400 gamma=32'd1;row=32'd281;
#400 gamma=32'd4;row=32'd529;
#400 gamma=32'd5;row=32'd289;
#400 gamma=32'd1;row=32'd143;
#400 gamma=32'd1;row=32'd201;
#400 gamma=32'd3;row=32'd509;
#400 gamma=32'd3;row=32'd380;
#400 gamma=32'd3;row=32'd39;
#400 gamma=32'd1;row=32'd372;
#400 gamma=32'd4;row=32'd196;
#400 gamma=32'd3;row=32'd547;
#400 gamma=32'd4;row=32'd94;
#400 gamma=32'd4;row=32'd486;
#400 gamma=32'd3;row=32'd288;
#400 gamma=32'd5;row=32'd64;
#400 gamma=32'd3;row=32'd355;
#400 gamma=32'd3;row=32'd529;
#400 gamma=32'd1;row=32'd521;
#400 gamma=32'd5;row=32'd92;
#400 gamma=32'd4;row=32'd62;
#400 gamma=32'd3;row=32'd362;
#400 gamma=32'd3;row=32'd383;
#400 gamma=32'd4;row=32'd458;
#400 gamma=32'd4;row=32'd434;
#400 gamma=32'd1;row=32'd187;
#400 gamma=32'd1;row=32'd391;
#400 gamma=32'd4;row=32'd37;
#400 gamma=32'd2;row=32'd433;
#400 gamma=32'd3;row=32'd6;
#400 gamma=32'd4;row=32'd165;
#400 gamma=32'd4;row=32'd436;
#400 gamma=32'd3;row=32'd48;
#400 gamma=32'd1;row=32'd162;
#400 gamma=32'd2;row=32'd59;
#400 gamma=32'd3;row=32'd247;
#400 gamma=32'd4;row=32'd180;
#400 gamma=32'd1;row=32'd552;
#400 gamma=32'd3;row=32'd84;
#400 gamma=32'd1;row=32'd224;
#400 gamma=32'd2;row=32'd209;
#400 gamma=32'd2;row=32'd487;
#400 gamma=32'd1;row=32'd440;
#400 gamma=32'd5;row=32'd357;
#400 gamma=32'd5;row=32'd472;
#400 gamma=32'd2;row=32'd129;
#400 gamma=32'd5;row=32'd276;
#400 gamma=32'd5;row=32'd190;
#400 gamma=32'd4;row=32'd47;
#400 gamma=32'd3;row=32'd487;
#400 gamma=32'd5;row=32'd17;
#400 gamma=32'd2;row=32'd291;
#400 gamma=32'd1;row=32'd3;
#400 gamma=32'd5;row=32'd236;
#400 gamma=32'd1;row=32'd544;
#400 gamma=32'd5;row=32'd340;
#400 gamma=32'd3;row=32'd80;
#400 gamma=32'd3;row=32'd88;
#400 gamma=32'd4;row=32'd92;
#400 gamma=32'd5;row=32'd435;
#400 gamma=32'd4;row=32'd430;
#400 gamma=32'd2;row=32'd345;
#400 gamma=32'd5;row=32'd509;
#400 gamma=32'd2;row=32'd304;
#400 gamma=32'd2;row=32'd163;
#400 gamma=32'd4;row=32'd205;
#400 gamma=32'd1;row=32'd383;
#400 gamma=32'd5;row=32'd179;
#400 gamma=32'd2;row=32'd549;
#400 gamma=32'd3;row=32'd426;
#400 gamma=32'd5;row=32'd208;
#400 gamma=32'd4;row=32'd427;
#400 gamma=32'd5;row=32'd257;
#400 gamma=32'd3;row=32'd407;
#400 gamma=32'd1;row=32'd461;
#400 gamma=32'd3;row=32'd307;
#400 gamma=32'd4;row=32'd302;
#400 gamma=32'd4;row=32'd80;
#400 gamma=32'd2;row=32'd502;
#400 gamma=32'd1;row=32'd287;
#400 gamma=32'd5;row=32'd531;
#400 gamma=32'd5;row=32'd54;
#400 gamma=32'd5;row=32'd195;
#400 gamma=32'd1;row=32'd275;
#400 gamma=32'd2;row=32'd207;
#400 gamma=32'd2;row=32'd514;
#400 gamma=32'd1;row=32'd243;
#400 gamma=32'd3;row=32'd517;
#400 gamma=32'd3;row=32'd176;
#400 gamma=32'd2;row=32'd380;
#400 gamma=32'd5;row=32'd42;
#400 gamma=32'd3;row=32'd431;
#400 gamma=32'd3;row=32'd231;
#400 gamma=32'd4;row=32'd553;
#400 gamma=32'd1;row=32'd100;
#400 gamma=32'd3;row=32'd237;
#400 gamma=32'd2;row=32'd77;
#400 gamma=32'd4;row=32'd493;
#400 gamma=32'd1;row=32'd296;
#400 gamma=32'd5;row=32'd251;
#400 gamma=32'd2;row=32'd516;
#400 gamma=32'd2;row=32'd323;
#400 gamma=32'd2;row=32'd292;
#400 gamma=32'd4;row=32'd140;
#400 gamma=32'd4;row=32'd328;
#400 gamma=32'd2;row=32'd495;
#400 gamma=32'd4;row=32'd315;
#400 gamma=32'd5;row=32'd370;
#400 gamma=32'd2;row=32'd292;
#400 gamma=32'd2;row=32'd278;
#400 gamma=32'd4;row=32'd210;
#400 gamma=32'd1;row=32'd507;
#400 gamma=32'd5;row=32'd417;
#400 gamma=32'd3;row=32'd100;
#400 gamma=32'd5;row=32'd73;
#400 gamma=32'd3;row=32'd157;
#400 gamma=32'd2;row=32'd225;
#400 gamma=32'd2;row=32'd194;
#400 gamma=32'd1;row=32'd152;
#400 gamma=32'd5;row=32'd40;
#400 gamma=32'd4;row=32'd373;
#400 gamma=32'd4;row=32'd244;
#400 gamma=32'd2;row=32'd135;
#400 gamma=32'd3;row=32'd49;
#400 gamma=32'd1;row=32'd94;
#400 gamma=32'd5;row=32'd47;
#400 gamma=32'd2;row=32'd558;
#400 gamma=32'd4;row=32'd444;
#400 gamma=32'd4;row=32'd280;
#400 gamma=32'd1;row=32'd296;
#400 gamma=32'd2;row=32'd13;
#400 gamma=32'd4;row=32'd264;
#400 gamma=32'd4;row=32'd15;
#400 gamma=32'd2;row=32'd253;
#400 gamma=32'd1;row=32'd195;
#400 gamma=32'd4;row=32'd211;
#400 gamma=32'd4;row=32'd130;
#400 gamma=32'd4;row=32'd233;
#400 gamma=32'd4;row=32'd448;
#400 gamma=32'd2;row=32'd352;
#400 gamma=32'd5;row=32'd320;
#400 gamma=32'd2;row=32'd96;
#400 gamma=32'd1;row=32'd226;
#400 gamma=32'd3;row=32'd21;
#400 gamma=32'd2;row=32'd26;
#400 gamma=32'd1;row=32'd128;
#400 gamma=32'd1;row=32'd459;
#400 gamma=32'd4;row=32'd115;
#400 gamma=32'd2;row=32'd192;
#400 gamma=32'd2;row=32'd158;
#400 gamma=32'd5;row=32'd463;
#400 gamma=32'd1;row=32'd121;
#400 gamma=32'd4;row=32'd97;
#400 gamma=32'd3;row=32'd57;
#400 gamma=32'd1;row=32'd282;
#400 gamma=32'd4;row=32'd414;
#400 gamma=32'd4;row=32'd126;
#400 gamma=32'd3;row=32'd380;
#400 gamma=32'd3;row=32'd296;
#400 gamma=32'd5;row=32'd267;
#400 gamma=32'd2;row=32'd74;
#400 gamma=32'd3;row=32'd273;
#400 gamma=32'd5;row=32'd41;
#400 gamma=32'd5;row=32'd319;
#400 gamma=32'd4;row=32'd476;
#400 gamma=32'd5;row=32'd504;
#400 gamma=32'd1;row=32'd196;
#400 gamma=32'd2;row=32'd457;
#400 gamma=32'd1;row=32'd393;
#400 gamma=32'd4;row=32'd15;
#400 gamma=32'd5;row=32'd31;
#400 gamma=32'd4;row=32'd118;
#400 gamma=32'd2;row=32'd453;
#400 gamma=32'd5;row=32'd223;
#400 gamma=32'd4;row=32'd205;
#400 gamma=32'd5;row=32'd73;
#400 gamma=32'd5;row=32'd534;
#400 gamma=32'd4;row=32'd50;
#400 gamma=32'd2;row=32'd358;
#400 gamma=32'd2;row=32'd81;
#400 gamma=32'd3;row=32'd192;
#400 gamma=32'd5;row=32'd372;
#400 gamma=32'd2;row=32'd96;
#400 gamma=32'd2;row=32'd169;
#400 gamma=32'd3;row=32'd517;
#400 gamma=32'd5;row=32'd120;
#400 gamma=32'd1;row=32'd370;
#400 gamma=32'd5;row=32'd117;
#400 gamma=32'd4;row=32'd431;
#400 gamma=32'd5;row=32'd232;
#400 gamma=32'd5;row=32'd19;
#400 gamma=32'd5;row=32'd392;
#400 gamma=32'd5;row=32'd379;
#400 gamma=32'd3;row=32'd90;
#400 gamma=32'd5;row=32'd537;
#400 gamma=32'd1;row=32'd334;
#400 gamma=32'd1;row=32'd479;
#400 gamma=32'd5;row=32'd462;
#400 gamma=32'd5;row=32'd0;
#400 gamma=32'd3;row=32'd415;
#400 gamma=32'd5;row=32'd39;
#400 gamma=32'd4;row=32'd12;
#400 gamma=32'd3;row=32'd316;
#400 gamma=32'd1;row=32'd508;
#400 gamma=32'd3;row=32'd209;
#400 gamma=32'd2;row=32'd254;
#400 gamma=32'd1;row=32'd180;
#400 gamma=32'd2;row=32'd327;
#400 gamma=32'd5;row=32'd434;
#400 gamma=32'd3;row=32'd179;
#400 gamma=32'd5;row=32'd163;
#400 gamma=32'd2;row=32'd309;
#400 gamma=32'd2;row=32'd203;
#400 gamma=32'd3;row=32'd415;
#400 gamma=32'd5;row=32'd520;
#400 gamma=32'd2;row=32'd9;
#400 gamma=32'd1;row=32'd394;
#400 gamma=32'd4;row=32'd438;
#400 gamma=32'd5;row=32'd300;
#400 gamma=32'd5;row=32'd123;
#400 gamma=32'd2;row=32'd410;
#400 gamma=32'd1;row=32'd48;
#400 gamma=32'd4;row=32'd147;
#400 gamma=32'd4;row=32'd340;
#400 gamma=32'd4;row=32'd364;
#400 gamma=32'd3;row=32'd251;
#400 gamma=32'd5;row=32'd256;
#400 gamma=32'd1;row=32'd233;
#400 gamma=32'd1;row=32'd180;
#400 gamma=32'd2;row=32'd95;
#400 gamma=32'd1;row=32'd512;
#400 gamma=32'd4;row=32'd4;
#400 gamma=32'd5;row=32'd249;
#400 gamma=32'd4;row=32'd265;
#400 gamma=32'd3;row=32'd359;
#400 gamma=32'd3;row=32'd212;
#400 gamma=32'd5;row=32'd352;
#400 gamma=32'd4;row=32'd342;
#400 gamma=32'd2;row=32'd360;
#400 gamma=32'd3;row=32'd444;
#400 gamma=32'd5;row=32'd469;
#400 gamma=32'd3;row=32'd171;
#400 gamma=32'd2;row=32'd216;
#400 gamma=32'd4;row=32'd42;
#400 gamma=32'd1;row=32'd545;
#400 gamma=32'd1;row=32'd111;
#400 gamma=32'd5;row=32'd441;
#400 gamma=32'd4;row=32'd66;
#400 gamma=32'd3;row=32'd232;
#400 gamma=32'd2;row=32'd300;
#400 gamma=32'd2;row=32'd529;
#400 gamma=32'd2;row=32'd243;
#400 gamma=32'd4;row=32'd333;
#400 gamma=32'd4;row=32'd402;
#400 gamma=32'd1;row=32'd542;
#400 gamma=32'd1;row=32'd59;
#400 gamma=32'd3;row=32'd299;
#400 gamma=32'd5;row=32'd552;
#400 gamma=32'd1;row=32'd109;
#400 gamma=32'd4;row=32'd555;
#400 gamma=32'd4;row=32'd81;
#400 gamma=32'd1;row=32'd482;
#400 gamma=32'd4;row=32'd34;
#400 gamma=32'd2;row=32'd550;
#400 gamma=32'd5;row=32'd163;
#400 gamma=32'd3;row=32'd458;
#400 gamma=32'd5;row=32'd299;
#400 gamma=32'd5;row=32'd224;
#400 gamma=32'd3;row=32'd208;
#400 gamma=32'd2;row=32'd263;
#400 gamma=32'd5;row=32'd53;
#400 gamma=32'd5;row=32'd374;
#400 gamma=32'd2;row=32'd553;
#400 gamma=32'd1;row=32'd58;
#400 gamma=32'd1;row=32'd544;
#400 gamma=32'd5;row=32'd263;
#400 gamma=32'd4;row=32'd349;
#400 gamma=32'd2;row=32'd192;
#400 gamma=32'd5;row=32'd276;
#400 gamma=32'd5;row=32'd128;
#400 gamma=32'd2;row=32'd126;
#400 gamma=32'd2;row=32'd376;
#400 gamma=32'd5;row=32'd325;
#400 gamma=32'd4;row=32'd309;
#400 gamma=32'd4;row=32'd556;
#400 gamma=32'd4;row=32'd187;
#400 gamma=32'd4;row=32'd291;
#400 gamma=32'd4;row=32'd485;
#400 gamma=32'd4;row=32'd275;
#400 gamma=32'd5;row=32'd55;
#400 gamma=32'd1;row=32'd477;
#400 gamma=32'd5;row=32'd290;
#400 gamma=32'd2;row=32'd475;
#400 gamma=32'd3;row=32'd280;
#400 gamma=32'd4;row=32'd393;
#400 gamma=32'd5;row=32'd461;
#400 gamma=32'd1;row=32'd182;
#400 gamma=32'd2;row=32'd308;
#400 gamma=32'd3;row=32'd215;
#400 gamma=32'd2;row=32'd105;
#400 gamma=32'd1;row=32'd36;
#400 gamma=32'd1;row=32'd355;
#400 gamma=32'd3;row=32'd191;
#400 gamma=32'd1;row=32'd81;
#400 gamma=32'd5;row=32'd454;
#400 gamma=32'd5;row=32'd540;
#400 gamma=32'd3;row=32'd269;
#400 gamma=32'd4;row=32'd139;
#400 gamma=32'd1;row=32'd157;
#400 gamma=32'd2;row=32'd181;
#400 gamma=32'd2;row=32'd160;
#400 gamma=32'd4;row=32'd401;
#400 gamma=32'd1;row=32'd152;
#400 gamma=32'd2;row=32'd62;
#400 gamma=32'd5;row=32'd464;
#400 gamma=32'd2;row=32'd453;
#400 gamma=32'd1;row=32'd137;
#400 gamma=32'd5;row=32'd49;
#400 gamma=32'd5;row=32'd265;
#400 gamma=32'd3;row=32'd431;
#400 gamma=32'd1;row=32'd243;
#400 gamma=32'd2;row=32'd506;
#400 gamma=32'd3;row=32'd404;
#400 gamma=32'd5;row=32'd112;
#400 gamma=32'd3;row=32'd375;
#400 gamma=32'd1;row=32'd556;
#400 gamma=32'd3;row=32'd45;
#400 gamma=32'd4;row=32'd95;
#400 gamma=32'd5;row=32'd151;
#400 gamma=32'd3;row=32'd16;
#400 gamma=32'd1;row=32'd142;
#400 gamma=32'd1;row=32'd506;
#400 gamma=32'd3;row=32'd536;
#400 gamma=32'd5;row=32'd538;
#400 gamma=32'd3;row=32'd82;
#400 gamma=32'd4;row=32'd280;
#400 gamma=32'd4;row=32'd505;
#400 gamma=32'd4;row=32'd69;
#400 gamma=32'd3;row=32'd338;
#400 gamma=32'd5;row=32'd474;
#400 gamma=32'd4;row=32'd68;
#400 gamma=32'd1;row=32'd69;
#400 gamma=32'd2;row=32'd7;
#400 gamma=32'd4;row=32'd268;
#400 gamma=32'd1;row=32'd535;
#400 gamma=32'd4;row=32'd41;
#400 gamma=32'd4;row=32'd534;
#400 gamma=32'd2;row=32'd472;
#400 gamma=32'd5;row=32'd70;
#400 gamma=32'd5;row=32'd150;
#400 gamma=32'd1;row=32'd172;
#400 gamma=32'd1;row=32'd143;
#400 gamma=32'd5;row=32'd529;
#400 gamma=32'd1;row=32'd541;
#400 gamma=32'd1;row=32'd426;
#400 gamma=32'd2;row=32'd319;
#400 gamma=32'd3;row=32'd172;
#400 gamma=32'd1;row=32'd80;
#400 gamma=32'd5;row=32'd400;
#400 gamma=32'd2;row=32'd524;
#400 gamma=32'd4;row=32'd199;
#400 gamma=32'd4;row=32'd52;
#400 gamma=32'd4;row=32'd80;
#400 gamma=32'd5;row=32'd195;
#400 gamma=32'd4;row=32'd516;
#400 gamma=32'd5;row=32'd490;
#400 gamma=32'd3;row=32'd135;
#400 gamma=32'd2;row=32'd12;
#400 gamma=32'd3;row=32'd542;
#400 gamma=32'd5;row=32'd177;
#400 gamma=32'd3;row=32'd427;
#400 gamma=32'd4;row=32'd500;
#400 gamma=32'd4;row=32'd207;
#400 gamma=32'd2;row=32'd223;
#400 gamma=32'd2;row=32'd299;
#400 gamma=32'd5;row=32'd6;
#400 gamma=32'd1;row=32'd382;
#400 gamma=32'd1;row=32'd260;
#400 gamma=32'd5;row=32'd491;
#400 gamma=32'd5;row=32'd295;
#400 gamma=32'd1;row=32'd485;
#400 gamma=32'd2;row=32'd540;
#400 gamma=32'd1;row=32'd479;
#400 gamma=32'd5;row=32'd357;
#400 gamma=32'd4;row=32'd145;
#400 gamma=32'd1;row=32'd348;
#400 gamma=32'd2;row=32'd525;
#400 gamma=32'd5;row=32'd187;
#400 gamma=32'd3;row=32'd418;
#400 gamma=32'd1;row=32'd200;
#400 gamma=32'd3;row=32'd167;
#400 gamma=32'd3;row=32'd245;
#400 gamma=32'd1;row=32'd197;
#400 gamma=32'd2;row=32'd61;
#400 gamma=32'd1;row=32'd527;
#400 gamma=32'd5;row=32'd272;
#400 gamma=32'd2;row=32'd408;
#400 gamma=32'd4;row=32'd40;
#400 gamma=32'd3;row=32'd376;
#400 gamma=32'd2;row=32'd188;
#400 gamma=32'd1;row=32'd481;
#400 gamma=32'd3;row=32'd205;
#400 gamma=32'd3;row=32'd457;
#400 gamma=32'd3;row=32'd441;
#400 gamma=32'd5;row=32'd26;
#400 gamma=32'd5;row=32'd133;
#400 gamma=32'd3;row=32'd303;
#400 gamma=32'd2;row=32'd233;
#400 gamma=32'd3;row=32'd77;
#400 gamma=32'd3;row=32'd109;
#400 gamma=32'd2;row=32'd47;
#400 gamma=32'd3;row=32'd170;
#400 gamma=32'd2;row=32'd35;
#400 gamma=32'd4;row=32'd183;
#400 gamma=32'd4;row=32'd310;
#400 gamma=32'd1;row=32'd490;
#400 gamma=32'd3;row=32'd37;
#400 gamma=32'd2;row=32'd198;
#400 gamma=32'd3;row=32'd266;
#400 gamma=32'd5;row=32'd137;
#400 gamma=32'd4;row=32'd127;
#400 gamma=32'd4;row=32'd479;
#400 gamma=32'd1;row=32'd171;
#400 gamma=32'd3;row=32'd474;
#400 gamma=32'd4;row=32'd330;
#400 gamma=32'd1;row=32'd470;
#400 gamma=32'd5;row=32'd77;
#400 gamma=32'd5;row=32'd81;
#400 gamma=32'd3;row=32'd285;
#400 gamma=32'd1;row=32'd294;
#400 gamma=32'd5;row=32'd546;
#400 gamma=32'd1;row=32'd379;
#400 gamma=32'd3;row=32'd536;
#400 gamma=32'd5;row=32'd374;
#400 gamma=32'd3;row=32'd140;
#400 gamma=32'd2;row=32'd376;
#400 gamma=32'd4;row=32'd39;
#400 gamma=32'd2;row=32'd55;
#400 gamma=32'd4;row=32'd20;
#400 gamma=32'd5;row=32'd554;
#400 gamma=32'd1;row=32'd86;
#400 gamma=32'd5;row=32'd44;
#400 gamma=32'd2;row=32'd201;
#400 gamma=32'd5;row=32'd125;
#400 gamma=32'd3;row=32'd510;
#400 gamma=32'd2;row=32'd417;
#400 gamma=32'd2;row=32'd81;
#400 gamma=32'd5;row=32'd26;
#400 gamma=32'd4;row=32'd377;
#400 gamma=32'd2;row=32'd87;
#400 gamma=32'd5;row=32'd382;
#400 gamma=32'd4;row=32'd525;
#400 gamma=32'd3;row=32'd329;
#400 gamma=32'd1;row=32'd549;
#400 gamma=32'd3;row=32'd176;
#400 gamma=32'd3;row=32'd1;
#400 gamma=32'd5;row=32'd256;
#400 gamma=32'd1;row=32'd110;
#400 gamma=32'd2;row=32'd526;
#400 gamma=32'd5;row=32'd532;
#400 gamma=32'd3;row=32'd102;
#400 gamma=32'd4;row=32'd510;
#400 gamma=32'd2;row=32'd355;
#400 gamma=32'd1;row=32'd38;
#400 gamma=32'd3;row=32'd199;
#400 gamma=32'd3;row=32'd100;
#400 gamma=32'd4;row=32'd454;
#400 gamma=32'd4;row=32'd298;
#400 gamma=32'd3;row=32'd182;
#400 gamma=32'd2;row=32'd300;
#400 gamma=32'd2;row=32'd133;
#400 gamma=32'd5;row=32'd485;
#400 gamma=32'd3;row=32'd275;
#400 gamma=32'd1;row=32'd352;
#400 gamma=32'd4;row=32'd82;
#400 gamma=32'd1;row=32'd248;
#400 gamma=32'd2;row=32'd36;
#400 gamma=32'd1;row=32'd108;
#400 gamma=32'd4;row=32'd376;
#400 gamma=32'd1;row=32'd303;
#400 gamma=32'd2;row=32'd518;
#400 gamma=32'd1;row=32'd532;
#400 gamma=32'd3;row=32'd462;
#400 gamma=32'd1;row=32'd514;
#400 gamma=32'd3;row=32'd396;
#400 gamma=32'd2;row=32'd435;
#400 gamma=32'd1;row=32'd456;
#400 gamma=32'd3;row=32'd201;
#400 gamma=32'd5;row=32'd496;
#400 gamma=32'd4;row=32'd104;
#400 gamma=32'd4;row=32'd543;
#400 gamma=32'd3;row=32'd126;
#400 gamma=32'd2;row=32'd493;
#400 gamma=32'd2;row=32'd198;
#400 gamma=32'd3;row=32'd124;
#400 gamma=32'd4;row=32'd11;
#400 gamma=32'd5;row=32'd396;
#400 gamma=32'd2;row=32'd335;
#400 gamma=32'd4;row=32'd87;
#400 gamma=32'd1;row=32'd144;
#400 gamma=32'd1;row=32'd310;
#400 gamma=32'd2;row=32'd408;
#400 gamma=32'd4;row=32'd174;
#400 gamma=32'd5;row=32'd6;
#400 gamma=32'd4;row=32'd236;
#400 gamma=32'd1;row=32'd286;
#400 gamma=32'd1;row=32'd269;
#400 gamma=32'd1;row=32'd484;
#400 gamma=32'd1;row=32'd294;
#400 gamma=32'd5;row=32'd22;
#400 gamma=32'd3;row=32'd189;
#400 gamma=32'd2;row=32'd72;
#400 gamma=32'd4;row=32'd301;
#400 gamma=32'd3;row=32'd431;
#400 gamma=32'd4;row=32'd368;
#400 gamma=32'd1;row=32'd76;
#400 gamma=32'd4;row=32'd460;
#400 gamma=32'd2;row=32'd44;
#400 gamma=32'd5;row=32'd24;
#400 gamma=32'd3;row=32'd23;
#400 gamma=32'd3;row=32'd12;
#400 gamma=32'd5;row=32'd536;
#400 gamma=32'd4;row=32'd344;
#400 gamma=32'd5;row=32'd553;
#400 gamma=32'd1;row=32'd113;
#400 gamma=32'd4;row=32'd13;
#400 gamma=32'd4;row=32'd166;
#400 gamma=32'd1;row=32'd402;
#400 gamma=32'd2;row=32'd347;
#400 gamma=32'd1;row=32'd27;
#400 gamma=32'd4;row=32'd208;
#400 gamma=32'd1;row=32'd439;
#400 gamma=32'd1;row=32'd482;
#400 gamma=32'd4;row=32'd341;
#400 gamma=32'd5;row=32'd77;
#400 gamma=32'd1;row=32'd257;
#400 gamma=32'd1;row=32'd461;
#400 gamma=32'd1;row=32'd41;
#400 gamma=32'd1;row=32'd532;
#400 gamma=32'd4;row=32'd502;
#400 gamma=32'd3;row=32'd136;
#400 gamma=32'd2;row=32'd394;
#400 gamma=32'd2;row=32'd302;
#400 gamma=32'd5;row=32'd372;
#400 gamma=32'd5;row=32'd117;
#400 gamma=32'd1;row=32'd428;
#400 gamma=32'd1;row=32'd424;
#400 gamma=32'd3;row=32'd482;
#400 gamma=32'd3;row=32'd515;
#400 gamma=32'd1;row=32'd303;
#400 gamma=32'd5;row=32'd231;
#400 gamma=32'd2;row=32'd36;
#400 gamma=32'd3;row=32'd48;
#400 gamma=32'd3;row=32'd18;
#400 gamma=32'd2;row=32'd505;
#400 gamma=32'd3;row=32'd160;
#400 gamma=32'd2;row=32'd350;
#400 gamma=32'd4;row=32'd160;
#400 gamma=32'd2;row=32'd427;
#400 gamma=32'd1;row=32'd417;
#400 gamma=32'd4;row=32'd272;
#400 gamma=32'd4;row=32'd441;
#400 gamma=32'd5;row=32'd163;
#400 gamma=32'd1;row=32'd50;
#400 gamma=32'd1;row=32'd549;
#400 gamma=32'd1;row=32'd224;
#400 gamma=32'd1;row=32'd193;
#400 gamma=32'd2;row=32'd120;
#400 gamma=32'd3;row=32'd305;
#400 gamma=32'd3;row=32'd227;
#400 gamma=32'd3;row=32'd250;
#400 gamma=32'd2;row=32'd302;
#400 gamma=32'd1;row=32'd50;
#400 gamma=32'd4;row=32'd345;
#400 gamma=32'd1;row=32'd41;
#400 gamma=32'd5;row=32'd149;
#400 gamma=32'd5;row=32'd80;
#400 gamma=32'd1;row=32'd222;
#400 gamma=32'd2;row=32'd540;
#400 gamma=32'd4;row=32'd327;
#400 gamma=32'd2;row=32'd300;
#400 gamma=32'd2;row=32'd479;
#400 gamma=32'd5;row=32'd217;
#400 gamma=32'd2;row=32'd520;
#400 gamma=32'd3;row=32'd524;
#400 gamma=32'd3;row=32'd300;
#400 gamma=32'd1;row=32'd33;
#400 gamma=32'd1;row=32'd497;
#400 gamma=32'd1;row=32'd83;
#400 gamma=32'd1;row=32'd35;
#400 gamma=32'd1;row=32'd474;
#400 gamma=32'd5;row=32'd28;
#400 gamma=32'd1;row=32'd52;
#400 gamma=32'd4;row=32'd287;
#400 gamma=32'd4;row=32'd137;
#400 gamma=32'd2;row=32'd77;
#400 gamma=32'd2;row=32'd521;
#400 gamma=32'd4;row=32'd57;
#400 gamma=32'd5;row=32'd111;
#400 gamma=32'd5;row=32'd314;
#400 gamma=32'd2;row=32'd283;
#400 gamma=32'd2;row=32'd408;
#400 gamma=32'd3;row=32'd75;
#400 gamma=32'd5;row=32'd497;
#400 gamma=32'd2;row=32'd148;
#400 gamma=32'd4;row=32'd411;
#400 gamma=32'd5;row=32'd420;
#400 gamma=32'd3;row=32'd271;
#400 gamma=32'd2;row=32'd525;
#400 gamma=32'd1;row=32'd467;
#400 gamma=32'd1;row=32'd102;
#400 gamma=32'd1;row=32'd489;
#400 gamma=32'd5;row=32'd382;
#400 gamma=32'd4;row=32'd142;
#400 gamma=32'd3;row=32'd506;
#400 gamma=32'd1;row=32'd169;
#400 gamma=32'd1;row=32'd72;
#400 gamma=32'd2;row=32'd430;
#400 gamma=32'd1;row=32'd46;
#400 gamma=32'd3;row=32'd43;
#400 gamma=32'd3;row=32'd284;
#400 gamma=32'd5;row=32'd281;
#400 gamma=32'd1;row=32'd39;
#400 gamma=32'd5;row=32'd366;
#400 gamma=32'd2;row=32'd263;
#400 gamma=32'd3;row=32'd284;
#400 gamma=32'd1;row=32'd527;
#400 gamma=32'd2;row=32'd8;
#400 gamma=32'd1;row=32'd309;
#400 gamma=32'd5;row=32'd246;
#400 gamma=32'd5;row=32'd119;
#400 gamma=32'd5;row=32'd510;
#400 gamma=32'd5;row=32'd373;
#400 gamma=32'd5;row=32'd451;
#400 gamma=32'd3;row=32'd105;
#400 gamma=32'd5;row=32'd96;
#400 gamma=32'd5;row=32'd407;
#400 gamma=32'd5;row=32'd527;
#400 gamma=32'd5;row=32'd501;
#400 gamma=32'd1;row=32'd549;
#400 gamma=32'd1;row=32'd156;
#400 gamma=32'd2;row=32'd388;
#400 gamma=32'd5;row=32'd283;
#400 gamma=32'd2;row=32'd321;
#400 gamma=32'd2;row=32'd474;
#400 gamma=32'd1;row=32'd46;
#400 gamma=32'd2;row=32'd390;
#400 gamma=32'd2;row=32'd206;
#400 gamma=32'd1;row=32'd131;
#400 gamma=32'd4;row=32'd501;
#400 gamma=32'd2;row=32'd226;
#400 gamma=32'd5;row=32'd65;
#400 gamma=32'd4;row=32'd449;
#400 gamma=32'd2;row=32'd389;
#400 gamma=32'd2;row=32'd7;
#400 gamma=32'd1;row=32'd14;
#400 gamma=32'd4;row=32'd61;
#400 gamma=32'd3;row=32'd71;
#400 gamma=32'd1;row=32'd136;
#400 gamma=32'd1;row=32'd501;
#400 gamma=32'd1;row=32'd166;
#400 gamma=32'd1;row=32'd213;
#400 gamma=32'd3;row=32'd63;
#400 gamma=32'd5;row=32'd424;
#400 gamma=32'd5;row=32'd215;
#400 gamma=32'd2;row=32'd412;
#400 gamma=32'd1;row=32'd463;
#400 gamma=32'd3;row=32'd417;
#400 gamma=32'd3;row=32'd4;
#400 gamma=32'd4;row=32'd177;
#400 gamma=32'd3;row=32'd542;
#400 gamma=32'd5;row=32'd346;
#400 gamma=32'd3;row=32'd442;
#400 gamma=32'd4;row=32'd357;
#400 gamma=32'd5;row=32'd290;
#400 gamma=32'd2;row=32'd206;
#400 gamma=32'd3;row=32'd401;
#400 gamma=32'd2;row=32'd307;
#400 gamma=32'd5;row=32'd123;
#400 gamma=32'd1;row=32'd510;
#400 gamma=32'd4;row=32'd537;
#400 gamma=32'd1;row=32'd239;
#400 gamma=32'd1;row=32'd88;
#400 gamma=32'd2;row=32'd549;
#400 gamma=32'd3;row=32'd54;
#400 gamma=32'd5;row=32'd187;
#400 gamma=32'd1;row=32'd244;
#400 gamma=32'd4;row=32'd494;
#400 gamma=32'd1;row=32'd97;
#400 gamma=32'd3;row=32'd7;
#400 gamma=32'd3;row=32'd267;
#400 gamma=32'd4;row=32'd361;
#400 gamma=32'd1;row=32'd210;
#400 gamma=32'd4;row=32'd393;
#400 gamma=32'd3;row=32'd264;
#400 gamma=32'd5;row=32'd511;
#400 gamma=32'd4;row=32'd435;
#400 gamma=32'd5;row=32'd253;
#400 gamma=32'd5;row=32'd468;
#400 gamma=32'd4;row=32'd335;
#400 gamma=32'd2;row=32'd49;
#400 gamma=32'd4;row=32'd436;
#400 gamma=32'd4;row=32'd538;
#400 gamma=32'd2;row=32'd177;
#400 gamma=32'd1;row=32'd39;
#400 gamma=32'd4;row=32'd79;
#400 gamma=32'd1;row=32'd60;
#400 gamma=32'd3;row=32'd119;
#400 gamma=32'd5;row=32'd72;
#400 gamma=32'd4;row=32'd269;
#400 gamma=32'd4;row=32'd16;
#400 gamma=32'd3;row=32'd199;
#400 gamma=32'd1;row=32'd429;
#400 gamma=32'd3;row=32'd40;
#400 gamma=32'd4;row=32'd330;
#400 gamma=32'd2;row=32'd341;
#400 gamma=32'd5;row=32'd194;
#400 gamma=32'd3;row=32'd476;
#400 gamma=32'd4;row=32'd23;
#400 gamma=32'd5;row=32'd408;
#400 gamma=32'd5;row=32'd285;
#400 gamma=32'd3;row=32'd4;
#400 gamma=32'd4;row=32'd193;
#400 gamma=32'd5;row=32'd509;
#400 gamma=32'd4;row=32'd119;
#400 gamma=32'd1;row=32'd204;
#400 gamma=32'd4;row=32'd143;
#400 gamma=32'd5;row=32'd198;
#400 gamma=32'd3;row=32'd202;
#400 gamma=32'd1;row=32'd104;
#400 gamma=32'd2;row=32'd100;
#400 gamma=32'd2;row=32'd530;
#400 gamma=32'd2;row=32'd55;
#400 gamma=32'd2;row=32'd209;
#400 gamma=32'd4;row=32'd193;
#400 gamma=32'd3;row=32'd300;
#400 gamma=32'd4;row=32'd191;
#400 gamma=32'd2;row=32'd385;
#400 gamma=32'd2;row=32'd357;
#400 gamma=32'd5;row=32'd70;
#400 gamma=32'd4;row=32'd444;
#400 gamma=32'd2;row=32'd200;
#400 gamma=32'd3;row=32'd359;
#400 gamma=32'd3;row=32'd463;
#400 gamma=32'd4;row=32'd494;
#400 gamma=32'd3;row=32'd532;
#400 gamma=32'd2;row=32'd331;
#400 gamma=32'd4;row=32'd326;
#400 gamma=32'd2;row=32'd35;
#400 gamma=32'd4;row=32'd115;
#400 gamma=32'd4;row=32'd314;
#400 gamma=32'd2;row=32'd237;
#400 gamma=32'd2;row=32'd272;
#400 gamma=32'd3;row=32'd465;
#400 gamma=32'd4;row=32'd37;
#400 gamma=32'd5;row=32'd475;
#400 gamma=32'd3;row=32'd328;
#400 gamma=32'd4;row=32'd267;
#400 gamma=32'd2;row=32'd196;
#400 gamma=32'd5;row=32'd372;
#400 gamma=32'd5;row=32'd214;
#400 gamma=32'd5;row=32'd376;
#400 gamma=32'd4;row=32'd163;
#400 gamma=32'd2;row=32'd490;
#400 gamma=32'd1;row=32'd83;
#400 gamma=32'd3;row=32'd207;
#400 gamma=32'd5;row=32'd289;
#400 gamma=32'd2;row=32'd75;
#400 gamma=32'd3;row=32'd123;
#400 gamma=32'd2;row=32'd292;
#400 gamma=32'd4;row=32'd369;
#400 gamma=32'd2;row=32'd509;
#400 gamma=32'd3;row=32'd366;
#400 gamma=32'd4;row=32'd26;
#400 gamma=32'd3;row=32'd158;
#400 gamma=32'd4;row=32'd551;
#400 gamma=32'd4;row=32'd458;
#400 gamma=32'd5;row=32'd536;
#400 gamma=32'd5;row=32'd227;
#400 gamma=32'd5;row=32'd398;
#400 gamma=32'd1;row=32'd432;
#400 gamma=32'd4;row=32'd453;
#400 gamma=32'd2;row=32'd310;
#400 gamma=32'd2;row=32'd257;
#400 gamma=32'd3;row=32'd105;
#400 gamma=32'd3;row=32'd212;
#400 gamma=32'd3;row=32'd293;
#400 gamma=32'd1;row=32'd41;
#400 gamma=32'd1;row=32'd533;
#400 gamma=32'd5;row=32'd247;
#400 gamma=32'd4;row=32'd50;
#400 gamma=32'd2;row=32'd83;
#400 gamma=32'd1;row=32'd427;
#400 gamma=32'd3;row=32'd433;
#400 gamma=32'd2;row=32'd509;
#400 gamma=32'd5;row=32'd461;
#400 gamma=32'd4;row=32'd402;
#400 gamma=32'd2;row=32'd351;
#400 gamma=32'd4;row=32'd194;
#400 gamma=32'd2;row=32'd362;
#400 gamma=32'd5;row=32'd341;
#400 gamma=32'd3;row=32'd513;
#400 gamma=32'd1;row=32'd226;
#400 gamma=32'd1;row=32'd104;
#400 gamma=32'd5;row=32'd219;
#400 gamma=32'd1;row=32'd552;
#400 gamma=32'd4;row=32'd44;
#400 gamma=32'd2;row=32'd423;
#400 gamma=32'd1;row=32'd17;
#400 gamma=32'd4;row=32'd281;
#400 gamma=32'd1;row=32'd369;
#400 gamma=32'd1;row=32'd196;
#400 gamma=32'd3;row=32'd310;
#400 gamma=32'd5;row=32'd96;
#400 gamma=32'd3;row=32'd62;
#400 gamma=32'd2;row=32'd247;
#400 gamma=32'd3;row=32'd551;
#400 gamma=32'd2;row=32'd30;
#400 gamma=32'd4;row=32'd397;
#400 gamma=32'd5;row=32'd24;
#400 gamma=32'd5;row=32'd36;
#400 gamma=32'd1;row=32'd354;
#400 gamma=32'd2;row=32'd273;
#400 gamma=32'd3;row=32'd123;
#400 gamma=32'd5;row=32'd394;
#400 gamma=32'd3;row=32'd517;
#400 gamma=32'd4;row=32'd415;
#400 gamma=32'd2;row=32'd58;
#400 gamma=32'd3;row=32'd429;
#400 gamma=32'd2;row=32'd245;
#400 gamma=32'd3;row=32'd273;
#400 gamma=32'd1;row=32'd381;
#400 gamma=32'd5;row=32'd67;
#400 gamma=32'd3;row=32'd17;
#400 gamma=32'd1;row=32'd91;
#400 gamma=32'd3;row=32'd188;
#400 gamma=32'd2;row=32'd354;
#400 gamma=32'd4;row=32'd13;
#400 gamma=32'd4;row=32'd329;
#400 gamma=32'd5;row=32'd172;
#400 gamma=32'd1;row=32'd323;
#400 gamma=32'd5;row=32'd466;
#400 gamma=32'd4;row=32'd441;
#400 gamma=32'd4;row=32'd9;
#400 gamma=32'd1;row=32'd310;
#400 gamma=32'd1;row=32'd134;
#400 gamma=32'd1;row=32'd283;
#400 gamma=32'd2;row=32'd106;
#400 gamma=32'd2;row=32'd120;
#400 gamma=32'd2;row=32'd525;
#400 gamma=32'd5;row=32'd445;
#400 gamma=32'd1;row=32'd144;
#400 gamma=32'd1;row=32'd258;
#400 gamma=32'd5;row=32'd245;
#400 gamma=32'd2;row=32'd559;
#400 gamma=32'd4;row=32'd184;
#400 gamma=32'd3;row=32'd310;
#400 gamma=32'd3;row=32'd358;
#400 gamma=32'd3;row=32'd353;
#400 gamma=32'd4;row=32'd309;
#400 gamma=32'd4;row=32'd401;
#400 gamma=32'd1;row=32'd471;
#400 gamma=32'd2;row=32'd331;
#400 gamma=32'd5;row=32'd281;
#400 gamma=32'd5;row=32'd14;
#400 gamma=32'd1;row=32'd186;
#400 gamma=32'd5;row=32'd206;
#400 gamma=32'd3;row=32'd162;
#400 gamma=32'd5;row=32'd360;
#400 gamma=32'd5;row=32'd510;
#400 gamma=32'd5;row=32'd518;
#400 gamma=32'd1;row=32'd385;
#400 gamma=32'd5;row=32'd431;
#400 gamma=32'd5;row=32'd429;
#400 gamma=32'd2;row=32'd526;
#400 gamma=32'd3;row=32'd385;
#400 gamma=32'd5;row=32'd345;
#400 gamma=32'd5;row=32'd403;
#400 gamma=32'd1;row=32'd477;
#400 gamma=32'd2;row=32'd150;
#400 gamma=32'd2;row=32'd120;
#400 gamma=32'd1;row=32'd454;
#400 gamma=32'd2;row=32'd217;
#400 gamma=32'd1;row=32'd150;
#400 gamma=32'd2;row=32'd483;
#400 gamma=32'd5;row=32'd66;
#400 gamma=32'd2;row=32'd553;
#400 gamma=32'd1;row=32'd538;
#400 gamma=32'd2;row=32'd19;
#400 gamma=32'd4;row=32'd529;
#400 gamma=32'd3;row=32'd157;
#400 gamma=32'd2;row=32'd551;
#400 gamma=32'd5;row=32'd2;
#400 gamma=32'd3;row=32'd108;
#400 gamma=32'd5;row=32'd490;
#400 gamma=32'd1;row=32'd413;
#400 gamma=32'd4;row=32'd269;
#400 gamma=32'd3;row=32'd490;
#400 gamma=32'd4;row=32'd304;
#400 gamma=32'd2;row=32'd18;
#400 gamma=32'd1;row=32'd495;
#400 gamma=32'd2;row=32'd194;
#400 gamma=32'd1;row=32'd492;
#400 gamma=32'd5;row=32'd336;
#400 gamma=32'd3;row=32'd442;
#400 gamma=32'd2;row=32'd312;
#400 gamma=32'd3;row=32'd72;
#400 gamma=32'd2;row=32'd276;
#400 gamma=32'd4;row=32'd304;
#400 gamma=32'd4;row=32'd114;
#400 gamma=32'd4;row=32'd414;
#400 gamma=32'd1;row=32'd179;
#400 gamma=32'd5;row=32'd418;
#400 gamma=32'd3;row=32'd48;
#400 gamma=32'd1;row=32'd151;
#400 gamma=32'd2;row=32'd111;
#400 gamma=32'd1;row=32'd17;
#400 gamma=32'd3;row=32'd237;
#400 gamma=32'd4;row=32'd84;
#400 gamma=32'd1;row=32'd216;
#400 gamma=32'd1;row=32'd208;
#400 gamma=32'd2;row=32'd415;
#400 gamma=32'd3;row=32'd359;
#400 gamma=32'd2;row=32'd141;
#400 gamma=32'd5;row=32'd534;
#400 gamma=32'd5;row=32'd198;
#400 gamma=32'd3;row=32'd96;
#400 gamma=32'd4;row=32'd326;
#400 gamma=32'd3;row=32'd130;
#400 gamma=32'd3;row=32'd209;
#400 gamma=32'd4;row=32'd246;
#400 gamma=32'd2;row=32'd524;
#400 gamma=32'd2;row=32'd388;
#400 gamma=32'd4;row=32'd369;
#400 gamma=32'd2;row=32'd10;
#400 gamma=32'd1;row=32'd86;
#400 gamma=32'd5;row=32'd240;
#400 gamma=32'd3;row=32'd319;
#400 gamma=32'd4;row=32'd329;
#400 gamma=32'd1;row=32'd86;
#400 gamma=32'd1;row=32'd376;
#400 gamma=32'd1;row=32'd8;
#400 gamma=32'd3;row=32'd251;
#400 gamma=32'd3;row=32'd21;
#400 gamma=32'd5;row=32'd444;
#400 gamma=32'd5;row=32'd537;
#400 gamma=32'd5;row=32'd359;
#400 gamma=32'd5;row=32'd192;
#400 gamma=32'd2;row=32'd55;
#400 gamma=32'd2;row=32'd453;
#400 gamma=32'd3;row=32'd251;
#400 gamma=32'd1;row=32'd207;
#400 gamma=32'd5;row=32'd557;
#400 gamma=32'd2;row=32'd275;
#400 gamma=32'd5;row=32'd24;
#400 gamma=32'd2;row=32'd276;
#400 gamma=32'd1;row=32'd118;
#400 gamma=32'd4;row=32'd329;
#400 gamma=32'd4;row=32'd407;
#400 gamma=32'd5;row=32'd15;
#400 gamma=32'd1;row=32'd95;
#400 gamma=32'd2;row=32'd379;
#400 gamma=32'd2;row=32'd62;
#400 gamma=32'd1;row=32'd552;
#400 gamma=32'd2;row=32'd61;
#400 gamma=32'd1;row=32'd128;
#400 gamma=32'd4;row=32'd114;
#400 gamma=32'd1;row=32'd191;
#400 gamma=32'd1;row=32'd309;
#400 gamma=32'd1;row=32'd380;
#400 gamma=32'd4;row=32'd336;
#400 gamma=32'd1;row=32'd463;
#400 gamma=32'd3;row=32'd549;
#400 gamma=32'd1;row=32'd92;
#400 gamma=32'd4;row=32'd538;
#400 gamma=32'd5;row=32'd208;
#400 gamma=32'd3;row=32'd237;
#400 gamma=32'd2;row=32'd117;
#400 gamma=32'd5;row=32'd165;
#400 gamma=32'd2;row=32'd342;
#400 gamma=32'd5;row=32'd407;
#400 gamma=32'd5;row=32'd313;
#400 gamma=32'd5;row=32'd116;
#400 gamma=32'd1;row=32'd310;
#400 gamma=32'd4;row=32'd383;
#400 gamma=32'd5;row=32'd57;
#400 gamma=32'd1;row=32'd214;
#400 gamma=32'd2;row=32'd131;
#400 gamma=32'd4;row=32'd305;
#400 gamma=32'd4;row=32'd363;
#400 gamma=32'd3;row=32'd512;
#400 gamma=32'd1;row=32'd325;
#400 gamma=32'd2;row=32'd513;
#400 gamma=32'd2;row=32'd509;
#400 gamma=32'd1;row=32'd446;
#400 gamma=32'd4;row=32'd539;
#400 gamma=32'd3;row=32'd82;
#400 gamma=32'd2;row=32'd275;
#400 gamma=32'd3;row=32'd225;
#400 gamma=32'd5;row=32'd428;
#400 gamma=32'd4;row=32'd91;
#400 gamma=32'd5;row=32'd325;
#400 gamma=32'd3;row=32'd46;
#400 gamma=32'd2;row=32'd30;
#400 gamma=32'd2;row=32'd207;
#400 gamma=32'd3;row=32'd558;
#400 gamma=32'd5;row=32'd74;
#400 gamma=32'd5;row=32'd299;
#400 gamma=32'd2;row=32'd85;
#400 gamma=32'd4;row=32'd71;
#400 gamma=32'd2;row=32'd9;
#400 gamma=32'd2;row=32'd235;
#400 gamma=32'd2;row=32'd260;
#400 gamma=32'd3;row=32'd427;
#400 gamma=32'd1;row=32'd48;
#400 gamma=32'd3;row=32'd466;
#400 gamma=32'd3;row=32'd418;
#400 gamma=32'd5;row=32'd514;
#400 gamma=32'd3;row=32'd30;
#400 gamma=32'd3;row=32'd252;
#400 gamma=32'd2;row=32'd408;
#400 gamma=32'd2;row=32'd150;
#400 gamma=32'd5;row=32'd209;
#400 gamma=32'd4;row=32'd488;
#400 gamma=32'd2;row=32'd395;
#400 gamma=32'd5;row=32'd142;
#400 gamma=32'd5;row=32'd329;
#400 gamma=32'd4;row=32'd511;
#400 gamma=32'd5;row=32'd462;
#400 gamma=32'd2;row=32'd14;
#400 gamma=32'd1;row=32'd195;
#400 gamma=32'd1;row=32'd84;
#400 gamma=32'd3;row=32'd212;
#400 gamma=32'd2;row=32'd40;
#400 gamma=32'd5;row=32'd18;
#400 gamma=32'd2;row=32'd499;
#400 gamma=32'd4;row=32'd157;
#400 gamma=32'd4;row=32'd435;
#400 gamma=32'd1;row=32'd112;
#400 gamma=32'd4;row=32'd164;
#400 gamma=32'd5;row=32'd472;
#400 gamma=32'd4;row=32'd385;
#400 gamma=32'd3;row=32'd373;
#400 gamma=32'd4;row=32'd20;
#400 gamma=32'd5;row=32'd246;
#400 gamma=32'd5;row=32'd68;
#400 gamma=32'd1;row=32'd56;
#400 gamma=32'd3;row=32'd472;
#400 gamma=32'd1;row=32'd498;
#400 gamma=32'd3;row=32'd347;
#400 gamma=32'd4;row=32'd230;
#400 gamma=32'd3;row=32'd440;
#400 gamma=32'd5;row=32'd59;
#400 gamma=32'd5;row=32'd264;
#400 gamma=32'd4;row=32'd427;
#400 gamma=32'd3;row=32'd84;
#400 gamma=32'd3;row=32'd314;
#400 gamma=32'd4;row=32'd480;
#400 gamma=32'd1;row=32'd100;
#400 gamma=32'd1;row=32'd26;
#400 gamma=32'd1;row=32'd31;
#400 gamma=32'd5;row=32'd544;
#400 gamma=32'd5;row=32'd338;
#400 gamma=32'd5;row=32'd109;
#400 gamma=32'd1;row=32'd27;
#400 gamma=32'd5;row=32'd26;
#400 gamma=32'd3;row=32'd142;
#400 gamma=32'd2;row=32'd513;
#400 gamma=32'd4;row=32'd355;
#400 gamma=32'd3;row=32'd537;
#400 gamma=32'd5;row=32'd453;
#400 gamma=32'd1;row=32'd203;
#400 gamma=32'd4;row=32'd336;
#400 gamma=32'd2;row=32'd118;
#400 gamma=32'd1;row=32'd332;
#400 gamma=32'd5;row=32'd400;
#400 gamma=32'd3;row=32'd196;
#400 gamma=32'd2;row=32'd92;
#400 gamma=32'd3;row=32'd174;
#400 gamma=32'd3;row=32'd515;
#400 gamma=32'd3;row=32'd495;
#400 gamma=32'd5;row=32'd333;
#400 gamma=32'd5;row=32'd91;
#400 gamma=32'd5;row=32'd290;
#400 gamma=32'd1;row=32'd493;
#400 gamma=32'd4;row=32'd277;
#400 gamma=32'd2;row=32'd223;
#400 gamma=32'd2;row=32'd1;
#400 gamma=32'd4;row=32'd73;
#400 gamma=32'd2;row=32'd75;
#400 gamma=32'd4;row=32'd16;
#400 gamma=32'd4;row=32'd340;
#400 gamma=32'd1;row=32'd315;
#400 gamma=32'd1;row=32'd444;
#400 gamma=32'd2;row=32'd152;
#400 gamma=32'd5;row=32'd340;
#400 gamma=32'd2;row=32'd396;
#400 gamma=32'd2;row=32'd414;
#400 gamma=32'd1;row=32'd100;
#400 gamma=32'd1;row=32'd300;
#400 gamma=32'd4;row=32'd316;
#400 gamma=32'd4;row=32'd220;
#400 gamma=32'd1;row=32'd165;
#400 gamma=32'd3;row=32'd209;
#400 gamma=32'd3;row=32'd285;
#400 gamma=32'd1;row=32'd197;
#400 gamma=32'd2;row=32'd232;
#400 gamma=32'd4;row=32'd4;
#400 gamma=32'd3;row=32'd2;
#400 gamma=32'd5;row=32'd102;
#400 gamma=32'd5;row=32'd469;
#400 gamma=32'd3;row=32'd185;
#400 gamma=32'd4;row=32'd32;
#400 gamma=32'd1;row=32'd384;
#400 gamma=32'd4;row=32'd547;
#400 gamma=32'd1;row=32'd402;
#400 gamma=32'd3;row=32'd115;
#400 gamma=32'd2;row=32'd552;
#400 gamma=32'd3;row=32'd362;
#400 gamma=32'd1;row=32'd446;
#400 gamma=32'd3;row=32'd479;
#400 gamma=32'd3;row=32'd410;
#400 gamma=32'd4;row=32'd544;
#400 gamma=32'd2;row=32'd103;
#400 gamma=32'd1;row=32'd464;
#400 gamma=32'd4;row=32'd519;
#400 gamma=32'd4;row=32'd51;
#400 gamma=32'd3;row=32'd393;
#400 gamma=32'd3;row=32'd506;
#400 gamma=32'd3;row=32'd199;
#400 gamma=32'd4;row=32'd373;
#400 gamma=32'd2;row=32'd95;
#400 gamma=32'd5;row=32'd338;
#400 gamma=32'd5;row=32'd415;
#400 gamma=32'd1;row=32'd531;
#400 gamma=32'd3;row=32'd490;
#400 gamma=32'd2;row=32'd254;
#400 gamma=32'd3;row=32'd250;
#400 gamma=32'd4;row=32'd541;
#400 gamma=32'd4;row=32'd40;
#400 gamma=32'd1;row=32'd123;
#400 gamma=32'd2;row=32'd247;
#400 gamma=32'd2;row=32'd494;
#400 gamma=32'd1;row=32'd129;
#400 gamma=32'd3;row=32'd185;
#400 gamma=32'd1;row=32'd119;
#400 gamma=32'd1;row=32'd237;
#400 gamma=32'd5;row=32'd448;
#400 gamma=32'd2;row=32'd159;
#400 gamma=32'd3;row=32'd519;
#400 gamma=32'd1;row=32'd538;
#400 gamma=32'd4;row=32'd153;
#400 gamma=32'd5;row=32'd210;
#400 gamma=32'd4;row=32'd468;
#400 gamma=32'd5;row=32'd535;
#400 gamma=32'd1;row=32'd47;
#400 gamma=32'd3;row=32'd128;
#400 gamma=32'd1;row=32'd461;
#400 gamma=32'd4;row=32'd228;
#400 gamma=32'd3;row=32'd226;
#400 gamma=32'd1;row=32'd526;
#400 gamma=32'd5;row=32'd127;
#400 gamma=32'd1;row=32'd557;
#400 gamma=32'd4;row=32'd6;
#400 gamma=32'd4;row=32'd76;
#400 gamma=32'd2;row=32'd474;
#400 gamma=32'd4;row=32'd234;
#400 gamma=32'd5;row=32'd276;
#400 gamma=32'd1;row=32'd340;
#400 gamma=32'd2;row=32'd113;
#400 gamma=32'd1;row=32'd102;
#400 gamma=32'd3;row=32'd393;
#400 gamma=32'd4;row=32'd279;
#400 gamma=32'd5;row=32'd438;
#400 gamma=32'd4;row=32'd179;
#400 gamma=32'd4;row=32'd122;
#400 gamma=32'd4;row=32'd368;
#400 gamma=32'd3;row=32'd14;
#400 gamma=32'd1;row=32'd201;
#400 gamma=32'd3;row=32'd301;
#400 gamma=32'd1;row=32'd458;
#400 gamma=32'd1;row=32'd173;
#400 gamma=32'd5;row=32'd552;
#400 gamma=32'd4;row=32'd38;
#400 gamma=32'd5;row=32'd498;
#400 gamma=32'd4;row=32'd399;
#400 gamma=32'd1;row=32'd265;
#400 gamma=32'd2;row=32'd305;
#400 gamma=32'd3;row=32'd455;
#400 gamma=32'd4;row=32'd37;
#400 gamma=32'd5;row=32'd7;
#400 gamma=32'd3;row=32'd240;
#400 gamma=32'd3;row=32'd461;
#400 gamma=32'd3;row=32'd138;
#400 gamma=32'd2;row=32'd95;
#400 gamma=32'd2;row=32'd177;
#400 gamma=32'd5;row=32'd264;
#400 gamma=32'd1;row=32'd530;
#400 gamma=32'd4;row=32'd310;
#400 gamma=32'd5;row=32'd1;
#400 gamma=32'd5;row=32'd93;
#400 gamma=32'd1;row=32'd469;
#400 gamma=32'd4;row=32'd465;
#400 gamma=32'd2;row=32'd274;
#400 gamma=32'd5;row=32'd310;
#400 gamma=32'd3;row=32'd363;
#400 gamma=32'd2;row=32'd396;
#400 gamma=32'd1;row=32'd551;
#400 gamma=32'd4;row=32'd488;
#400 gamma=32'd3;row=32'd174;
#400 gamma=32'd1;row=32'd253;
#400 gamma=32'd4;row=32'd275;
#400 gamma=32'd2;row=32'd4;
#400 gamma=32'd1;row=32'd277;
#400 gamma=32'd1;row=32'd521;
#400 gamma=32'd2;row=32'd486;
#400 gamma=32'd2;row=32'd213;
#400 gamma=32'd5;row=32'd310;
#400 gamma=32'd1;row=32'd174;
#400 gamma=32'd4;row=32'd112;
#400 gamma=32'd3;row=32'd220;
#400 gamma=32'd3;row=32'd98;
#400 gamma=32'd5;row=32'd337;
#400 gamma=32'd5;row=32'd288;
#400 gamma=32'd4;row=32'd223;
#400 gamma=32'd5;row=32'd377;
#400 gamma=32'd2;row=32'd345;
#400 gamma=32'd3;row=32'd366;
#400 gamma=32'd3;row=32'd246;
#400 gamma=32'd2;row=32'd35;
#400 gamma=32'd4;row=32'd31;
#400 gamma=32'd3;row=32'd418;
#400 gamma=32'd5;row=32'd239;
#400 gamma=32'd4;row=32'd248;
#400 gamma=32'd3;row=32'd296;
#400 gamma=32'd4;row=32'd495;
#400 gamma=32'd4;row=32'd558;
#400 gamma=32'd1;row=32'd442;
#400 gamma=32'd4;row=32'd7;
#400 gamma=32'd1;row=32'd128;
#400 gamma=32'd1;row=32'd339;
#400 gamma=32'd2;row=32'd81;
#400 gamma=32'd2;row=32'd187;
#400 gamma=32'd5;row=32'd518;
#400 gamma=32'd5;row=32'd191;
#400 gamma=32'd2;row=32'd438;
#400 gamma=32'd4;row=32'd173;
#400 gamma=32'd4;row=32'd179;
#400 gamma=32'd4;row=32'd89;
#400 gamma=32'd4;row=32'd526;
#400 gamma=32'd3;row=32'd278;
#400 gamma=32'd3;row=32'd454;
#400 gamma=32'd4;row=32'd68;
#400 gamma=32'd1;row=32'd231;
#400 gamma=32'd5;row=32'd453;
#400 gamma=32'd4;row=32'd447;
#400 gamma=32'd3;row=32'd195;
// dense
#800 gamma=1;row=1;
#800 gamma=1;row=1; 
#7600 gamma=1; row=1;
end





endmodule
